`ifdef _SPD_TB_MATCH
module spd_tb_decoder (
// input
phy_mode_bit, gen, refclk_fsel, ref_clk_ring_sel, reg_fbck_sel,
ring_dis,
// output
pll_rate_sel_tx_expected, tx_ck_sel_lane_expected,
tx_vddcal_rate_en_lane_expected, tx_speed_div_lane_expected,
tx_reg_speed_trk_clk_lane_expected, tx_reg_speed_trk_data_lane_expected,
tx_em_ctrl_reg_en_lane_expected, tx_em_ctrl_pipe_sel_lane_expected,
tx_em_pre_en_lane_expected, tx_em_pre_ctrl_lane_expected,
tx_em_po_en_lane_expected, tx_em_po_ctrl_lane_expected,
slewrate_en_lane_expected, slewctrl1_lane_expected,
slewctrl0_lane_expected, tx_train_pat_sel_lane_expected,
train_pat_num_lane_expected, tx_train_pat_toggle_lane_expected,
packet_sync_dis_lane_expected, sync_det_dis_lane_expected,
pll_rate_sel_rx_expected, rx_ck_sel_lane_expected,
rx_vddcal_rate_en_lane_expected, rx_speed_div_lane_expected,
dtl_clk_speedup_lane_expected, intpi_lane_expected,
intpr_lane_expected, dll_freq_sel_lane_expected, eom_dll_freq_sel_lane_expected,
align90_8g_en_lane_expected, rx_reg0p9_speed_track_clk_lane_expected,
rx_reg0p9_speed_track_clk_half_lane_expected, rx_reg0p9_speed_track_data_lane_expected,
rx_selmufi_lane_expected, rx_selmuff_lane_expected,
reg_selmupi_lane_expected, reg_selmupf_lane_expected,
rx_rxclk_25m_ctrl_lane_expected, rx_rxclk_25m_div1p5_en_lane_expected,
rx_rxclk_25m_div_lane_expected, rx_rxclk_25m_fix_div_en_lane_expected,
dtl_clk_mode_lane_expected, rx_foffset_extra_m_lane_expected,
init_rxfoffs_lane_expected, pu_f1p_d_e_lane_expected,
pu_f1n_d_e_lane_expected, pu_f1p_s_e_lane_expected,
pu_f1n_s_e_lane_expected, pu_f1p_d_o_lane_expected,
pu_f1n_d_o_lane_expected, pu_f1p_s_o_lane_expected,
pu_f1n_s_o_lane_expected, path_disable_edge_lane_expected,
dfe_f1_pol_en_d_lane_expected, dfe_f1_pol_en_s_lane_expected,
dfe_f1_pol_d_lane_expected, dfe_f1_pol_s_lane_expected,
reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected, reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected,
reg_ana_rx_dfe_f1_pol_d_force_lane_expected, reg_ana_rx_dfe_f1_pol_s_force_lane_expected,
reg_dfe_full_rate_mode_lane_expected, reg_dfe_dis_lane_expected,
reg_dfe_tap_settle_scale_lane_expected, ffe_data_rate_lane_expected,
ffe_res1_sel_lane_expected, ffe_cap1_sel_lane_expected,
ffe_res2_sel_e_lane_expected, ffe_res2_sel_o_lane_expected,
ffe_cap2_sel_e_lane_expected, ffe_cap2_sel_o_lane_expected,
rxdll_temp_a_lane_expected, rxdll_temp_b_lane_expected,
pll_reg_sel_expected, pll_rate_sel_expected, fbdiv_expected,
fbdiv_cal_expected, refdiv_expected, vind_band_sel_expected,
div_1g_expected, div_1g_fbck_expected, icp_lc_expected,
pll_lpfr_expected, pll_lpfc_expected, intpi_lcpll_expected,
tx_intpr_expected, init_txfoffs_expected, speed_thresh_expected,
lccap_usb_expected, ssc_acc_factor_expected, ssc_step_125ppm_expected,
ssc_m_expected, ref_clk_ring_sel_expected, clk1g_refclk_sel_expected,
pll_refdiv_ring_expected, pll_fbdiv_ring_expected,
pll_fbdiv_ring_fbck_expected, icp_ring_expected, pll_speed_thresh_ring_expected,
fbdiv_cal_ring_expected, intpi_ring_expected, tx_intpr_ring_expected,
pll_band_sel_ring_expected, pll_lpf_c1_sel_ring_expected,
pll_lpf_c2_sel_ring_expected, pll_lpf_r1_sel_ring_expected,
init_txfoffs_ring_expected, init_txfoffs_ring_fbck_expected,
ssc_acc_factor_ring_expected, ssc_step_125ppm_ring_expected,
ssc_m_ring_expected
);

// parameters
parameter SATA = 3'd0;
parameter SAS = 3'd1;
parameter FC = 3'd2;
parameter PCIE = 3'd3;
parameter SERDES = 3'd4;
parameter USB = 3'd5;


input         [2:0]     phy_mode_bit;
input         [3:0]     gen;
input         [4:0]     refclk_fsel;
input                   ref_clk_ring_sel;
input                   reg_fbck_sel;
input                   ring_dis;

output        [3 : 0]   pll_rate_sel_tx_expected;
output                  tx_ck_sel_lane_expected;
output                  tx_vddcal_rate_en_lane_expected;
output        [2 : 0]   tx_speed_div_lane_expected;
output        [2 : 0]   tx_reg_speed_trk_clk_lane_expected;
output        [2 : 0]   tx_reg_speed_trk_data_lane_expected;
output                  tx_em_ctrl_reg_en_lane_expected;
output                  tx_em_ctrl_pipe_sel_lane_expected;
output                  tx_em_pre_en_lane_expected;
output        [3 : 0]   tx_em_pre_ctrl_lane_expected;
output                  tx_em_po_en_lane_expected;
output        [3 : 0]   tx_em_po_ctrl_lane_expected;
output        [1 : 0]   slewrate_en_lane_expected;
output        [1 : 0]   slewctrl1_lane_expected;
output        [1 : 0]   slewctrl0_lane_expected;
output        [1 : 0]   tx_train_pat_sel_lane_expected;
output        [8 : 0]   train_pat_num_lane_expected;
output                  tx_train_pat_toggle_lane_expected;
output                  packet_sync_dis_lane_expected;
output                  sync_det_dis_lane_expected;
output        [3 : 0]   pll_rate_sel_rx_expected;
output                  rx_ck_sel_lane_expected;
output                  rx_vddcal_rate_en_lane_expected;
output        [2 : 0]   rx_speed_div_lane_expected;
output        [2 : 0]   dtl_clk_speedup_lane_expected;
output        [3 : 0]   intpi_lane_expected;
output        [1 : 0]   intpr_lane_expected;
output        [2 : 0]   dll_freq_sel_lane_expected;
output        [2 : 0]   eom_dll_freq_sel_lane_expected;
output                  align90_8g_en_lane_expected;
output        [2 : 0]   rx_reg0p9_speed_track_clk_lane_expected;
output                  rx_reg0p9_speed_track_clk_half_lane_expected;
output        [2 : 0]   rx_reg0p9_speed_track_data_lane_expected;
output        [2 : 0]   rx_selmufi_lane_expected;
output        [2 : 0]   rx_selmuff_lane_expected;
output        [3 : 0]   reg_selmupi_lane_expected;
output        [3 : 0]   reg_selmupf_lane_expected;
output        [1 : 0]   rx_rxclk_25m_ctrl_lane_expected;
output                  rx_rxclk_25m_div1p5_en_lane_expected;
output        [7 : 0]   rx_rxclk_25m_div_lane_expected;
output                  rx_rxclk_25m_fix_div_en_lane_expected;
output        [1 : 0]   dtl_clk_mode_lane_expected;
output        [13 : 0]  rx_foffset_extra_m_lane_expected;
output        [9 : 0]   init_rxfoffs_lane_expected;
output                  pu_f1p_d_e_lane_expected;
output                  pu_f1n_d_e_lane_expected;
output                  pu_f1p_s_e_lane_expected;
output                  pu_f1n_s_e_lane_expected;
output                  pu_f1p_d_o_lane_expected;
output                  pu_f1n_d_o_lane_expected;
output                  pu_f1p_s_o_lane_expected;
output                  pu_f1n_s_o_lane_expected;
output                  path_disable_edge_lane_expected;
output                  dfe_f1_pol_en_d_lane_expected;
output                  dfe_f1_pol_en_s_lane_expected;
output                  dfe_f1_pol_d_lane_expected;
output                  dfe_f1_pol_s_lane_expected;
output                  reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected;
output                  reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected;
output                  reg_ana_rx_dfe_f1_pol_d_force_lane_expected;
output                  reg_ana_rx_dfe_f1_pol_s_force_lane_expected;
output                  reg_dfe_full_rate_mode_lane_expected;
output                  reg_dfe_dis_lane_expected;
output        [1 : 0]   reg_dfe_tap_settle_scale_lane_expected;
output        [3 : 0]   ffe_data_rate_lane_expected;
output        [3 : 0]   ffe_res1_sel_lane_expected;
output        [3 : 0]   ffe_cap1_sel_lane_expected;
output        [3 : 0]   ffe_res2_sel_e_lane_expected;
output        [3 : 0]   ffe_res2_sel_o_lane_expected;
output        [3 : 0]   ffe_cap2_sel_e_lane_expected;
output        [3 : 0]   ffe_cap2_sel_o_lane_expected;
output        [7 : 0]   rxdll_temp_a_lane_expected;
output        [7 : 0]   rxdll_temp_b_lane_expected;
output        [2 : 0]   pll_reg_sel_expected;
output        [3 : 0]   pll_rate_sel_expected;
output        [9 : 0]   fbdiv_expected;
output        [9 : 0]   fbdiv_cal_expected;
output        [3 : 0]   refdiv_expected;
output                  vind_band_sel_expected;
output        [9 : 0]   div_1g_expected;
output        [9 : 0]   div_1g_fbck_expected;
output        [4 : 0]   icp_lc_expected;
output        [1 : 0]   pll_lpfr_expected;
output        [1 : 0]   pll_lpfc_expected;
output        [3 : 0]   intpi_lcpll_expected;
output        [1 : 0]   tx_intpr_expected;
output        [9 : 0]   init_txfoffs_expected;
output        [11 : 0]  speed_thresh_expected;
output                  lccap_usb_expected;
output                  ssc_acc_factor_expected;
output        [3 : 0]   ssc_step_125ppm_expected;
output        [12 : 0]  ssc_m_expected;
output                  ref_clk_ring_sel_expected;
output                  clk1g_refclk_sel_expected;
output        [3 : 0]   pll_refdiv_ring_expected;
output        [9 : 0]   pll_fbdiv_ring_expected;
output        [9 : 0]   pll_fbdiv_ring_fbck_expected;
output        [3 : 0]   icp_ring_expected;
output        [8 : 0]   pll_speed_thresh_ring_expected;
output        [9 : 0]   fbdiv_cal_ring_expected;
output        [3 : 0]   intpi_ring_expected;
output        [1 : 0]   tx_intpr_ring_expected;
output                  pll_band_sel_ring_expected;
output        [1 : 0]   pll_lpf_c1_sel_ring_expected;
output        [1 : 0]   pll_lpf_c2_sel_ring_expected;
output        [2 : 0]   pll_lpf_r1_sel_ring_expected;
output        [9 : 0]   init_txfoffs_ring_expected;
output        [9 : 0]   init_txfoffs_ring_fbck_expected;
output                  ssc_acc_factor_ring_expected;
output        [3 : 0]   ssc_step_125ppm_ring_expected;
output        [12 : 0]  ssc_m_ring_expected;

wire          [4:0]     refclk_fsel_ring;

assign refclk_fsel_ring = (ref_clk_ring_sel == 1'b1) ? refclk_fsel : 5'd8;


reg           [3 : 0]   pll_rate_sel_tx_expected;
reg                     tx_ck_sel_lane_expected;
reg                     tx_vddcal_rate_en_lane_expected;
reg           [2 : 0]   tx_speed_div_lane_expected;
reg           [2 : 0]   tx_reg_speed_trk_clk_lane_expected;
reg           [2 : 0]   tx_reg_speed_trk_data_lane_expected;
reg                     tx_em_ctrl_reg_en_lane_expected;
reg                     tx_em_ctrl_pipe_sel_lane_expected;
reg                     tx_em_pre_en_lane_expected;
reg           [3 : 0]   tx_em_pre_ctrl_lane_expected;
reg                     tx_em_po_en_lane_expected;
reg           [3 : 0]   tx_em_po_ctrl_lane_expected;
reg           [1 : 0]   slewrate_en_lane_expected;
reg           [1 : 0]   slewctrl1_lane_expected;
reg           [1 : 0]   slewctrl0_lane_expected;
reg           [1 : 0]   tx_train_pat_sel_lane_expected;
reg           [8 : 0]   train_pat_num_lane_expected;
reg                     tx_train_pat_toggle_lane_expected;
reg                     packet_sync_dis_lane_expected;
reg                     sync_det_dis_lane_expected;
reg           [3 : 0]   pll_rate_sel_rx_expected;
reg                     rx_ck_sel_lane_expected;
reg                     rx_vddcal_rate_en_lane_expected;
reg           [2 : 0]   rx_speed_div_lane_expected;
reg           [2 : 0]   dtl_clk_speedup_lane_expected;
reg           [3 : 0]   intpi_lane_expected;
reg           [1 : 0]   intpr_lane_expected;
reg           [2 : 0]   dll_freq_sel_lane_expected;
reg           [2 : 0]   eom_dll_freq_sel_lane_expected;
reg                     align90_8g_en_lane_expected;
reg           [2 : 0]   rx_reg0p9_speed_track_clk_lane_expected;
reg                     rx_reg0p9_speed_track_clk_half_lane_expected;
reg           [2 : 0]   rx_reg0p9_speed_track_data_lane_expected;
reg           [2 : 0]   rx_selmufi_lane_expected;
reg           [2 : 0]   rx_selmuff_lane_expected;
reg           [3 : 0]   reg_selmupi_lane_expected;
reg           [3 : 0]   reg_selmupf_lane_expected;
reg           [1 : 0]   rx_rxclk_25m_ctrl_lane_expected;
reg                     rx_rxclk_25m_div1p5_en_lane_expected;
reg           [7 : 0]   rx_rxclk_25m_div_lane_expected;
reg                     rx_rxclk_25m_fix_div_en_lane_expected;
reg           [1 : 0]   dtl_clk_mode_lane_expected;
reg           [13 : 0]  rx_foffset_extra_m_lane_expected;
reg           [9 : 0]   init_rxfoffs_lane_expected;
reg                     pu_f1p_d_e_lane_expected;
reg                     pu_f1n_d_e_lane_expected;
reg                     pu_f1p_s_e_lane_expected;
reg                     pu_f1n_s_e_lane_expected;
reg                     pu_f1p_d_o_lane_expected;
reg                     pu_f1n_d_o_lane_expected;
reg                     pu_f1p_s_o_lane_expected;
reg                     pu_f1n_s_o_lane_expected;
reg                     path_disable_edge_lane_expected;
reg                     dfe_f1_pol_en_d_lane_expected;
reg                     dfe_f1_pol_en_s_lane_expected;
reg                     dfe_f1_pol_d_lane_expected;
reg                     dfe_f1_pol_s_lane_expected;
reg                     reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected;
reg                     reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected;
reg                     reg_ana_rx_dfe_f1_pol_d_force_lane_expected;
reg                     reg_ana_rx_dfe_f1_pol_s_force_lane_expected;
reg                     reg_dfe_full_rate_mode_lane_expected;
reg                     reg_dfe_dis_lane_expected;
reg           [1 : 0]   reg_dfe_tap_settle_scale_lane_expected;
reg           [3 : 0]   ffe_data_rate_lane_expected;
reg           [3 : 0]   ffe_res1_sel_lane_expected;
reg           [3 : 0]   ffe_cap1_sel_lane_expected;
reg           [3 : 0]   ffe_res2_sel_e_lane_expected;
reg           [3 : 0]   ffe_res2_sel_o_lane_expected;
reg           [3 : 0]   ffe_cap2_sel_e_lane_expected;
reg           [3 : 0]   ffe_cap2_sel_o_lane_expected;
reg           [7 : 0]   rxdll_temp_a_lane_expected;
reg           [7 : 0]   rxdll_temp_b_lane_expected;
reg           [2 : 0]   pll_reg_sel_expected;
reg           [3 : 0]   pll_rate_sel_expected;
reg           [9 : 0]   fbdiv_expected;
reg           [9 : 0]   fbdiv_cal_expected;
reg           [3 : 0]   refdiv_expected;
reg                     vind_band_sel_expected;
reg           [9 : 0]   div_1g_expected;
reg           [9 : 0]   div_1g_fbck_expected;
reg           [4 : 0]   icp_lc_expected;
reg           [1 : 0]   pll_lpfr_expected;
reg           [1 : 0]   pll_lpfc_expected;
reg           [3 : 0]   intpi_lcpll_expected;
reg           [1 : 0]   tx_intpr_expected;
reg           [9 : 0]   init_txfoffs_expected;
reg           [11 : 0]  speed_thresh_expected;
reg                     lccap_usb_expected;
reg                     ssc_acc_factor_expected;
reg           [3 : 0]   ssc_step_125ppm_expected;
reg           [12 : 0]  ssc_m_expected;
reg                     ref_clk_ring_sel_expected;
reg                     clk1g_refclk_sel_expected;
reg           [3 : 0]   pll_refdiv_ring_expected;
reg           [9 : 0]   pll_fbdiv_ring_expected;
reg           [9 : 0]   pll_fbdiv_ring_fbck_expected;
reg           [3 : 0]   icp_ring_expected;
reg           [8 : 0]   pll_speed_thresh_ring_expected;
reg           [9 : 0]   fbdiv_cal_ring_expected;
reg           [3 : 0]   intpi_ring_expected;
reg           [1 : 0]   tx_intpr_ring_expected;
reg                     pll_band_sel_ring_expected;
reg           [1 : 0]   pll_lpf_c1_sel_ring_expected;
reg           [1 : 0]   pll_lpf_c2_sel_ring_expected;
reg           [2 : 0]   pll_lpf_r1_sel_ring_expected;
reg           [9 : 0]   init_txfoffs_ring_expected;
reg           [9 : 0]   init_txfoffs_ring_fbck_expected;
reg                     ssc_acc_factor_ring_expected;
reg           [3 : 0]   ssc_step_125ppm_ring_expected;
reg           [12 : 0]  ssc_m_ring_expected;

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : pll_rate_sel_tx_expected = 4'b0000;
  {USB, 4'd2} : pll_rate_sel_tx_expected = 4'b0000;
  {SERDES, 4'd0} : pll_rate_sel_tx_expected = 4'b0000;
  {SERDES, 4'd1} : pll_rate_sel_tx_expected = 4'b0011;
  {SERDES, 4'd2} : pll_rate_sel_tx_expected = 4'b0001;
  {SERDES, 4'd3} : pll_rate_sel_tx_expected = 4'b0011;
  {SERDES, 4'd4} : pll_rate_sel_tx_expected = 4'b0001;
  {SERDES, 4'd5} : pll_rate_sel_tx_expected = 4'b0010;
  {SERDES, 4'd6} : pll_rate_sel_tx_expected = 4'b0011;
  {SERDES, 4'd7} : pll_rate_sel_tx_expected = 4'b0100;
  {SERDES, 4'd8} : pll_rate_sel_tx_expected = 4'b0101;
  {SERDES, 4'd9} : pll_rate_sel_tx_expected = 4'b0110;
  {SERDES, 4'd12} : pll_rate_sel_tx_expected = 4'b0000;
  {SERDES, 4'd13} : pll_rate_sel_tx_expected = 4'b0001;
  {SAS, 4'd0} : pll_rate_sel_tx_expected = 4'b0001;
  {SAS, 4'd1} : pll_rate_sel_tx_expected = 4'b0001;
  {SAS, 4'd2} : pll_rate_sel_tx_expected = 4'b0001;
  {SAS, 4'd3} : pll_rate_sel_tx_expected = 4'b0001;
  {SAS, 4'd4} : pll_rate_sel_tx_expected = 4'b0000;
  {PCIE, 4'd0} : pll_rate_sel_tx_expected = 4'b0001;
  {PCIE, 4'd1} : pll_rate_sel_tx_expected = 4'b0001;
  {PCIE, 4'd2} : pll_rate_sel_tx_expected = 4'b0000;
  {PCIE, 4'd3} : pll_rate_sel_tx_expected = 4'b0000;
default: pll_rate_sel_tx_expected = 4'bzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : tx_ck_sel_lane_expected = 1'b0;
  {USB, 4'd2} : tx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd0} : tx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd1} : tx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd2} : tx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd3} : tx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd4} : tx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd5} : tx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd6} : tx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd7} : tx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd8} : tx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd9} : tx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd12} : tx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd13} : tx_ck_sel_lane_expected = 1'b0;
  {SAS, 4'd0} : tx_ck_sel_lane_expected = 1'b0;
  {SAS, 4'd1} : tx_ck_sel_lane_expected = 1'b0;
  {SAS, 4'd2} : tx_ck_sel_lane_expected = 1'b0;
  {SAS, 4'd3} : tx_ck_sel_lane_expected = 1'b0;
  {SAS, 4'd4} : tx_ck_sel_lane_expected = 1'b0;
  {PCIE, 4'd0} : tx_ck_sel_lane_expected = 1'b1;
  {PCIE, 4'd1} : tx_ck_sel_lane_expected = 1'b1;
  {PCIE, 4'd2} : tx_ck_sel_lane_expected = 1'b0;
  {PCIE, 4'd3} : tx_ck_sel_lane_expected = 1'b0;
default: tx_ck_sel_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : tx_vddcal_rate_en_lane_expected = 1'b1;
  {USB, 4'd2} : tx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd0} : tx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd1} : tx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd2} : tx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd3} : tx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd4} : tx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd5} : tx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd6} : tx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd7} : tx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd8} : tx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd9} : tx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd12} : tx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd13} : tx_vddcal_rate_en_lane_expected = 1'b1;
  {SAS, 4'd0} : tx_vddcal_rate_en_lane_expected = 1'b1;
  {SAS, 4'd1} : tx_vddcal_rate_en_lane_expected = 1'b1;
  {SAS, 4'd2} : tx_vddcal_rate_en_lane_expected = 1'b1;
  {SAS, 4'd3} : tx_vddcal_rate_en_lane_expected = 1'b1;
  {SAS, 4'd4} : tx_vddcal_rate_en_lane_expected = 1'b1;
  {PCIE, 4'd0} : tx_vddcal_rate_en_lane_expected = 1'b1;
  {PCIE, 4'd1} : tx_vddcal_rate_en_lane_expected = 1'b1;
  {PCIE, 4'd2} : tx_vddcal_rate_en_lane_expected = 1'b1;
  {PCIE, 4'd3} : tx_vddcal_rate_en_lane_expected = 1'b1;
default: tx_vddcal_rate_en_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : tx_speed_div_lane_expected = 3'b010;
  {USB, 4'd2} : tx_speed_div_lane_expected = 3'b001;
  {SERDES, 4'd0} : tx_speed_div_lane_expected = 3'b100;
  {SERDES, 4'd1} : tx_speed_div_lane_expected = 3'b011;
  {SERDES, 4'd2} : tx_speed_div_lane_expected = 3'b010;
  {SERDES, 4'd3} : tx_speed_div_lane_expected = 3'b010;
  {SERDES, 4'd4} : tx_speed_div_lane_expected = 3'b001;
  {SERDES, 4'd5} : tx_speed_div_lane_expected = 3'b001;
  {SERDES, 4'd6} : tx_speed_div_lane_expected = 3'b001;
  {SERDES, 4'd7} : tx_speed_div_lane_expected = 3'b000;
  {SERDES, 4'd8} : tx_speed_div_lane_expected = 3'b000;
  {SERDES, 4'd9} : tx_speed_div_lane_expected = 3'b000;
  {SERDES, 4'd12} : tx_speed_div_lane_expected = 3'b011;
  {SERDES, 4'd13} : tx_speed_div_lane_expected = 3'b000;
  {SAS, 4'd0} : tx_speed_div_lane_expected = 3'b100;
  {SAS, 4'd1} : tx_speed_div_lane_expected = 3'b011;
  {SAS, 4'd2} : tx_speed_div_lane_expected = 3'b010;
  {SAS, 4'd3} : tx_speed_div_lane_expected = 3'b001;
  {SAS, 4'd4} : tx_speed_div_lane_expected = 3'b000;
  {PCIE, 4'd0} : tx_speed_div_lane_expected = 3'b011;
  {PCIE, 4'd1} : tx_speed_div_lane_expected = 3'b010;
  {PCIE, 4'd2} : tx_speed_div_lane_expected = 3'b001;
  {PCIE, 4'd3} : tx_speed_div_lane_expected = 3'b000;
default: tx_speed_div_lane_expected = 3'bzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : tx_reg_speed_trk_clk_lane_expected = 3'b011;
  {USB, 4'd2} : tx_reg_speed_trk_clk_lane_expected = 3'b011;
  {SERDES, 4'd0} : tx_reg_speed_trk_clk_lane_expected = 3'b001;
  {SERDES, 4'd1} : tx_reg_speed_trk_clk_lane_expected = 3'b001;
  {SERDES, 4'd2} : tx_reg_speed_trk_clk_lane_expected = 3'b011;
  {SERDES, 4'd3} : tx_reg_speed_trk_clk_lane_expected = 3'b001;
  {SERDES, 4'd4} : tx_reg_speed_trk_clk_lane_expected = 3'b011;
  {SERDES, 4'd5} : tx_reg_speed_trk_clk_lane_expected = 3'b011;
  {SERDES, 4'd6} : tx_reg_speed_trk_clk_lane_expected = 3'b011;
  {SERDES, 4'd7} : tx_reg_speed_trk_clk_lane_expected = 3'b111;
  {SERDES, 4'd8} : tx_reg_speed_trk_clk_lane_expected = 3'b111;
  {SERDES, 4'd9} : tx_reg_speed_trk_clk_lane_expected = 3'b111;
  {SERDES, 4'd12} : tx_reg_speed_trk_clk_lane_expected = 3'b011;
  {SERDES, 4'd13} : tx_reg_speed_trk_clk_lane_expected = 3'b110;
  {SAS, 4'd0} : tx_reg_speed_trk_clk_lane_expected = 3'b001;
  {SAS, 4'd1} : tx_reg_speed_trk_clk_lane_expected = 3'b001;
  {SAS, 4'd2} : tx_reg_speed_trk_clk_lane_expected = 3'b001;
  {SAS, 4'd3} : tx_reg_speed_trk_clk_lane_expected = 3'b011;
  {SAS, 4'd4} : tx_reg_speed_trk_clk_lane_expected = 3'b110;
  {PCIE, 4'd0} : tx_reg_speed_trk_clk_lane_expected = 3'b011;
  {PCIE, 4'd1} : tx_reg_speed_trk_clk_lane_expected = 3'b011;
  {PCIE, 4'd2} : tx_reg_speed_trk_clk_lane_expected = 3'b010;
  {PCIE, 4'd3} : tx_reg_speed_trk_clk_lane_expected = 3'b100;
default: tx_reg_speed_trk_clk_lane_expected = 3'bzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : tx_reg_speed_trk_data_lane_expected = 3'b011;
  {USB, 4'd2} : tx_reg_speed_trk_data_lane_expected = 3'b011;
  {SERDES, 4'd0} : tx_reg_speed_trk_data_lane_expected = 3'b001;
  {SERDES, 4'd1} : tx_reg_speed_trk_data_lane_expected = 3'b001;
  {SERDES, 4'd2} : tx_reg_speed_trk_data_lane_expected = 3'b011;
  {SERDES, 4'd3} : tx_reg_speed_trk_data_lane_expected = 3'b001;
  {SERDES, 4'd4} : tx_reg_speed_trk_data_lane_expected = 3'b011;
  {SERDES, 4'd5} : tx_reg_speed_trk_data_lane_expected = 3'b011;
  {SERDES, 4'd6} : tx_reg_speed_trk_data_lane_expected = 3'b011;
  {SERDES, 4'd7} : tx_reg_speed_trk_data_lane_expected = 3'b111;
  {SERDES, 4'd8} : tx_reg_speed_trk_data_lane_expected = 3'b111;
  {SERDES, 4'd9} : tx_reg_speed_trk_data_lane_expected = 3'b111;
  {SERDES, 4'd12} : tx_reg_speed_trk_data_lane_expected = 3'b011;
  {SERDES, 4'd13} : tx_reg_speed_trk_data_lane_expected = 3'b110;
  {SAS, 4'd0} : tx_reg_speed_trk_data_lane_expected = 3'b001;
  {SAS, 4'd1} : tx_reg_speed_trk_data_lane_expected = 3'b001;
  {SAS, 4'd2} : tx_reg_speed_trk_data_lane_expected = 3'b001;
  {SAS, 4'd3} : tx_reg_speed_trk_data_lane_expected = 3'b011;
  {SAS, 4'd4} : tx_reg_speed_trk_data_lane_expected = 3'b110;
  {PCIE, 4'd0} : tx_reg_speed_trk_data_lane_expected = 3'b011;
  {PCIE, 4'd1} : tx_reg_speed_trk_data_lane_expected = 3'b011;
  {PCIE, 4'd2} : tx_reg_speed_trk_data_lane_expected = 3'b010;
  {PCIE, 4'd3} : tx_reg_speed_trk_data_lane_expected = 3'b100;
default: tx_reg_speed_trk_data_lane_expected = 3'bzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : tx_em_ctrl_reg_en_lane_expected = 1'b0;
  {USB, 4'd2} : tx_em_ctrl_reg_en_lane_expected = 1'b0;
  {SERDES, 4'd0} : tx_em_ctrl_reg_en_lane_expected = 1'b1;
  {SERDES, 4'd1} : tx_em_ctrl_reg_en_lane_expected = 1'b1;
  {SERDES, 4'd2} : tx_em_ctrl_reg_en_lane_expected = 1'b0;
  {SERDES, 4'd3} : tx_em_ctrl_reg_en_lane_expected = 1'b1;
  {SERDES, 4'd4} : tx_em_ctrl_reg_en_lane_expected = 1'b1;
  {SERDES, 4'd5} : tx_em_ctrl_reg_en_lane_expected = 1'b1;
  {SERDES, 4'd6} : tx_em_ctrl_reg_en_lane_expected = 1'b1;
  {SERDES, 4'd7} : tx_em_ctrl_reg_en_lane_expected = 1'b1;
  {SERDES, 4'd8} : tx_em_ctrl_reg_en_lane_expected = 1'b1;
  {SERDES, 4'd9} : tx_em_ctrl_reg_en_lane_expected = 1'b1;
  {SERDES, 4'd12} : tx_em_ctrl_reg_en_lane_expected = 1'b0;
  {SERDES, 4'd13} : tx_em_ctrl_reg_en_lane_expected = 1'b1;
  {SAS, 4'd0} : tx_em_ctrl_reg_en_lane_expected = 1'b1;
  {SAS, 4'd1} : tx_em_ctrl_reg_en_lane_expected = 1'b1;
  {SAS, 4'd2} : tx_em_ctrl_reg_en_lane_expected = 1'b1;
  {SAS, 4'd3} : tx_em_ctrl_reg_en_lane_expected = 1'b1;
  {SAS, 4'd4} : tx_em_ctrl_reg_en_lane_expected = 1'b1;
  {PCIE, 4'd0} : tx_em_ctrl_reg_en_lane_expected = 1'b0;
  {PCIE, 4'd1} : tx_em_ctrl_reg_en_lane_expected = 1'b0;
  {PCIE, 4'd2} : tx_em_ctrl_reg_en_lane_expected = 1'b0;
  {PCIE, 4'd3} : tx_em_ctrl_reg_en_lane_expected = 1'b0;
default: tx_em_ctrl_reg_en_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : tx_em_ctrl_pipe_sel_lane_expected = 1'b0;
  {USB, 4'd2} : tx_em_ctrl_pipe_sel_lane_expected = 1'b0;
  {SERDES, 4'd0} : tx_em_ctrl_pipe_sel_lane_expected = 1'b0;
  {SERDES, 4'd1} : tx_em_ctrl_pipe_sel_lane_expected = 1'b0;
  {SERDES, 4'd2} : tx_em_ctrl_pipe_sel_lane_expected = 1'b0;
  {SERDES, 4'd3} : tx_em_ctrl_pipe_sel_lane_expected = 1'b0;
  {SERDES, 4'd4} : tx_em_ctrl_pipe_sel_lane_expected = 1'b0;
  {SERDES, 4'd5} : tx_em_ctrl_pipe_sel_lane_expected = 1'b0;
  {SERDES, 4'd6} : tx_em_ctrl_pipe_sel_lane_expected = 1'b0;
  {SERDES, 4'd7} : tx_em_ctrl_pipe_sel_lane_expected = 1'b0;
  {SERDES, 4'd8} : tx_em_ctrl_pipe_sel_lane_expected = 1'b0;
  {SERDES, 4'd9} : tx_em_ctrl_pipe_sel_lane_expected = 1'b0;
  {SERDES, 4'd12} : tx_em_ctrl_pipe_sel_lane_expected = 1'b0;
  {SERDES, 4'd13} : tx_em_ctrl_pipe_sel_lane_expected = 1'b0;
  {SAS, 4'd0} : tx_em_ctrl_pipe_sel_lane_expected = 1'b0;
  {SAS, 4'd1} : tx_em_ctrl_pipe_sel_lane_expected = 1'b0;
  {SAS, 4'd2} : tx_em_ctrl_pipe_sel_lane_expected = 1'b0;
  {SAS, 4'd3} : tx_em_ctrl_pipe_sel_lane_expected = 1'b0;
  {SAS, 4'd4} : tx_em_ctrl_pipe_sel_lane_expected = 1'b0;
  {PCIE, 4'd0} : tx_em_ctrl_pipe_sel_lane_expected = 1'b0;
  {PCIE, 4'd1} : tx_em_ctrl_pipe_sel_lane_expected = 1'b0;
  {PCIE, 4'd2} : tx_em_ctrl_pipe_sel_lane_expected = 1'b1;
  {PCIE, 4'd3} : tx_em_ctrl_pipe_sel_lane_expected = 1'b1;
default: tx_em_ctrl_pipe_sel_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : tx_em_pre_en_lane_expected = 1'b0;
  {USB, 4'd2} : tx_em_pre_en_lane_expected = 1'b0;
  {SERDES, 4'd0} : tx_em_pre_en_lane_expected = 1'b0;
  {SERDES, 4'd1} : tx_em_pre_en_lane_expected = 1'b0;
  {SERDES, 4'd2} : tx_em_pre_en_lane_expected = 1'b1;
  {SERDES, 4'd3} : tx_em_pre_en_lane_expected = 1'b1;
  {SERDES, 4'd4} : tx_em_pre_en_lane_expected = 1'b1;
  {SERDES, 4'd5} : tx_em_pre_en_lane_expected = 1'b1;
  {SERDES, 4'd6} : tx_em_pre_en_lane_expected = 1'b1;
  {SERDES, 4'd7} : tx_em_pre_en_lane_expected = 1'b1;
  {SERDES, 4'd8} : tx_em_pre_en_lane_expected = 1'b1;
  {SERDES, 4'd9} : tx_em_pre_en_lane_expected = 1'b1;
  {SERDES, 4'd12} : tx_em_pre_en_lane_expected = 1'b0;
  {SERDES, 4'd13} : tx_em_pre_en_lane_expected = 1'b1;
  {SAS, 4'd0} : tx_em_pre_en_lane_expected = 1'b0;
  {SAS, 4'd1} : tx_em_pre_en_lane_expected = 1'b0;
  {SAS, 4'd2} : tx_em_pre_en_lane_expected = 1'b0;
  {SAS, 4'd3} : tx_em_pre_en_lane_expected = 1'b1;
  {SAS, 4'd4} : tx_em_pre_en_lane_expected = 1'b1;
  {PCIE, 4'd0} : tx_em_pre_en_lane_expected = 1'b0;
  {PCIE, 4'd1} : tx_em_pre_en_lane_expected = 1'b0;
  {PCIE, 4'd2} : tx_em_pre_en_lane_expected = 1'b1;
  {PCIE, 4'd3} : tx_em_pre_en_lane_expected = 1'b1;
default: tx_em_pre_en_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : tx_em_pre_ctrl_lane_expected = 4'b1111;
  {USB, 4'd2} : tx_em_pre_ctrl_lane_expected = 4'b1111;
  {SERDES, 4'd0} : tx_em_pre_ctrl_lane_expected = 4'b1111;
  {SERDES, 4'd1} : tx_em_pre_ctrl_lane_expected = 4'b1011;
  {SERDES, 4'd2} : tx_em_pre_ctrl_lane_expected = 4'b0000;
  {SERDES, 4'd3} : tx_em_pre_ctrl_lane_expected = 4'b0000;
  {SERDES, 4'd4} : tx_em_pre_ctrl_lane_expected = 4'b0000;
  {SERDES, 4'd5} : tx_em_pre_ctrl_lane_expected = 4'b0000;
  {SERDES, 4'd6} : tx_em_pre_ctrl_lane_expected = 4'b0000;
  {SERDES, 4'd7} : tx_em_pre_ctrl_lane_expected = 4'b0000;
  {SERDES, 4'd8} : tx_em_pre_ctrl_lane_expected = 4'b0000;
  {SERDES, 4'd9} : tx_em_pre_ctrl_lane_expected = 4'b0000;
  {SERDES, 4'd12} : tx_em_pre_ctrl_lane_expected = 4'b1000;
  {SERDES, 4'd13} : tx_em_pre_ctrl_lane_expected = 4'b0000;
  {SAS, 4'd0} : tx_em_pre_ctrl_lane_expected = 4'b1000;
  {SAS, 4'd1} : tx_em_pre_ctrl_lane_expected = 4'b1011;
  {SAS, 4'd2} : tx_em_pre_ctrl_lane_expected = 4'b1011;
  {SAS, 4'd3} : tx_em_pre_ctrl_lane_expected = 4'b0000;
  {SAS, 4'd4} : tx_em_pre_ctrl_lane_expected = 4'b0000;
  {PCIE, 4'd0} : tx_em_pre_ctrl_lane_expected = 4'b1000;
  {PCIE, 4'd1} : tx_em_pre_ctrl_lane_expected = 4'b1011;
  {PCIE, 4'd2} : tx_em_pre_ctrl_lane_expected = 4'b0000;
  {PCIE, 4'd3} : tx_em_pre_ctrl_lane_expected = 4'b0000;
default: tx_em_pre_ctrl_lane_expected = 4'bzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : tx_em_po_en_lane_expected = 1'b0;
  {USB, 4'd2} : tx_em_po_en_lane_expected = 1'b0;
  {SERDES, 4'd0} : tx_em_po_en_lane_expected = 1'b0;
  {SERDES, 4'd1} : tx_em_po_en_lane_expected = 1'b0;
  {SERDES, 4'd2} : tx_em_po_en_lane_expected = 1'b1;
  {SERDES, 4'd3} : tx_em_po_en_lane_expected = 1'b1;
  {SERDES, 4'd4} : tx_em_po_en_lane_expected = 1'b1;
  {SERDES, 4'd5} : tx_em_po_en_lane_expected = 1'b1;
  {SERDES, 4'd6} : tx_em_po_en_lane_expected = 1'b1;
  {SERDES, 4'd7} : tx_em_po_en_lane_expected = 1'b1;
  {SERDES, 4'd8} : tx_em_po_en_lane_expected = 1'b1;
  {SERDES, 4'd9} : tx_em_po_en_lane_expected = 1'b1;
  {SERDES, 4'd12} : tx_em_po_en_lane_expected = 1'b0;
  {SERDES, 4'd13} : tx_em_po_en_lane_expected = 1'b1;
  {SAS, 4'd0} : tx_em_po_en_lane_expected = 1'b0;
  {SAS, 4'd1} : tx_em_po_en_lane_expected = 1'b0;
  {SAS, 4'd2} : tx_em_po_en_lane_expected = 1'b0;
  {SAS, 4'd3} : tx_em_po_en_lane_expected = 1'b1;
  {SAS, 4'd4} : tx_em_po_en_lane_expected = 1'b1;
  {PCIE, 4'd0} : tx_em_po_en_lane_expected = 1'b0;
  {PCIE, 4'd1} : tx_em_po_en_lane_expected = 1'b0;
  {PCIE, 4'd2} : tx_em_po_en_lane_expected = 1'b1;
  {PCIE, 4'd3} : tx_em_po_en_lane_expected = 1'b1;
default: tx_em_po_en_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : tx_em_po_ctrl_lane_expected = 4'b1111;
  {USB, 4'd2} : tx_em_po_ctrl_lane_expected = 4'b1111;
  {SERDES, 4'd0} : tx_em_po_ctrl_lane_expected = 4'b1111;
  {SERDES, 4'd1} : tx_em_po_ctrl_lane_expected = 4'b1111;
  {SERDES, 4'd2} : tx_em_po_ctrl_lane_expected = 4'b0000;
  {SERDES, 4'd3} : tx_em_po_ctrl_lane_expected = 4'b0000;
  {SERDES, 4'd4} : tx_em_po_ctrl_lane_expected = 4'b0000;
  {SERDES, 4'd5} : tx_em_po_ctrl_lane_expected = 4'b0000;
  {SERDES, 4'd6} : tx_em_po_ctrl_lane_expected = 4'b0000;
  {SERDES, 4'd7} : tx_em_po_ctrl_lane_expected = 4'b0000;
  {SERDES, 4'd8} : tx_em_po_ctrl_lane_expected = 4'b0000;
  {SERDES, 4'd9} : tx_em_po_ctrl_lane_expected = 4'b0000;
  {SERDES, 4'd12} : tx_em_po_ctrl_lane_expected = 4'b1111;
  {SERDES, 4'd13} : tx_em_po_ctrl_lane_expected = 4'b0000;
  {SAS, 4'd0} : tx_em_po_ctrl_lane_expected = 4'b1111;
  {SAS, 4'd1} : tx_em_po_ctrl_lane_expected = 4'b1111;
  {SAS, 4'd2} : tx_em_po_ctrl_lane_expected = 4'b1111;
  {SAS, 4'd3} : tx_em_po_ctrl_lane_expected = 4'b0000;
  {SAS, 4'd4} : tx_em_po_ctrl_lane_expected = 4'b0000;
  {PCIE, 4'd0} : tx_em_po_ctrl_lane_expected = 4'b1111;
  {PCIE, 4'd1} : tx_em_po_ctrl_lane_expected = 4'b1111;
  {PCIE, 4'd2} : tx_em_po_ctrl_lane_expected = 4'b0000;
  {PCIE, 4'd3} : tx_em_po_ctrl_lane_expected = 4'b0000;
default: tx_em_po_ctrl_lane_expected = 4'bzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : slewrate_en_lane_expected = 2'b00;
  {USB, 4'd2} : slewrate_en_lane_expected = 2'b00;
  {SERDES, 4'd0} : slewrate_en_lane_expected = 2'b00;
  {SERDES, 4'd1} : slewrate_en_lane_expected = 2'b11;
  {SERDES, 4'd2} : slewrate_en_lane_expected = 2'b11;
  {SERDES, 4'd3} : slewrate_en_lane_expected = 2'b11;
  {SERDES, 4'd4} : slewrate_en_lane_expected = 2'b00;
  {SERDES, 4'd5} : slewrate_en_lane_expected = 2'b01;
  {SERDES, 4'd6} : slewrate_en_lane_expected = 2'b00;
  {SERDES, 4'd7} : slewrate_en_lane_expected = 2'b00;
  {SERDES, 4'd8} : slewrate_en_lane_expected = 2'b00;
  {SERDES, 4'd9} : slewrate_en_lane_expected = 2'b00;
  {SERDES, 4'd12} : slewrate_en_lane_expected = 2'b11;
  {SERDES, 4'd13} : slewrate_en_lane_expected = 2'b00;
  {SAS, 4'd0} : slewrate_en_lane_expected = 2'b11;
  {SAS, 4'd1} : slewrate_en_lane_expected = 2'b11;
  {SAS, 4'd2} : slewrate_en_lane_expected = 2'b11;
  {SAS, 4'd3} : slewrate_en_lane_expected = 2'b00;
  {SAS, 4'd4} : slewrate_en_lane_expected = 2'b00;
  {PCIE, 4'd0} : slewrate_en_lane_expected = 2'b11;
  {PCIE, 4'd1} : slewrate_en_lane_expected = 2'b11;
  {PCIE, 4'd2} : slewrate_en_lane_expected = 2'b00;
  {PCIE, 4'd3} : slewrate_en_lane_expected = 2'b00;
default: slewrate_en_lane_expected = 2'bzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : slewctrl1_lane_expected = 2'b00;
  {USB, 4'd2} : slewctrl1_lane_expected = 2'b00;
  {SERDES, 4'd0} : slewctrl1_lane_expected = 2'b00;
  {SERDES, 4'd1} : slewctrl1_lane_expected = 2'b10;
  {SERDES, 4'd2} : slewctrl1_lane_expected = 2'b10;
  {SERDES, 4'd3} : slewctrl1_lane_expected = 2'b10;
  {SERDES, 4'd4} : slewctrl1_lane_expected = 2'b00;
  {SERDES, 4'd5} : slewctrl1_lane_expected = 2'b00;
  {SERDES, 4'd6} : slewctrl1_lane_expected = 2'b00;
  {SERDES, 4'd7} : slewctrl1_lane_expected = 2'b00;
  {SERDES, 4'd8} : slewctrl1_lane_expected = 2'b00;
  {SERDES, 4'd9} : slewctrl1_lane_expected = 2'b00;
  {SERDES, 4'd12} : slewctrl1_lane_expected = 2'b10;
  {SERDES, 4'd13} : slewctrl1_lane_expected = 2'b00;
  {SAS, 4'd0} : slewctrl1_lane_expected = 2'b10;
  {SAS, 4'd1} : slewctrl1_lane_expected = 2'b10;
  {SAS, 4'd2} : slewctrl1_lane_expected = 2'b10;
  {SAS, 4'd3} : slewctrl1_lane_expected = 2'b00;
  {SAS, 4'd4} : slewctrl1_lane_expected = 2'b00;
  {PCIE, 4'd0} : slewctrl1_lane_expected = 2'b10;
  {PCIE, 4'd1} : slewctrl1_lane_expected = 2'b10;
  {PCIE, 4'd2} : slewctrl1_lane_expected = 2'b00;
  {PCIE, 4'd3} : slewctrl1_lane_expected = 2'b00;
default: slewctrl1_lane_expected = 2'bzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : slewctrl0_lane_expected = 2'b00;
  {USB, 4'd2} : slewctrl0_lane_expected = 2'b00;
  {SERDES, 4'd0} : slewctrl0_lane_expected = 2'b00;
  {SERDES, 4'd1} : slewctrl0_lane_expected = 2'b01;
  {SERDES, 4'd2} : slewctrl0_lane_expected = 2'b01;
  {SERDES, 4'd3} : slewctrl0_lane_expected = 2'b01;
  {SERDES, 4'd4} : slewctrl0_lane_expected = 2'b00;
  {SERDES, 4'd5} : slewctrl0_lane_expected = 2'b00;
  {SERDES, 4'd6} : slewctrl0_lane_expected = 2'b00;
  {SERDES, 4'd7} : slewctrl0_lane_expected = 2'b00;
  {SERDES, 4'd8} : slewctrl0_lane_expected = 2'b00;
  {SERDES, 4'd9} : slewctrl0_lane_expected = 2'b00;
  {SERDES, 4'd12} : slewctrl0_lane_expected = 2'b01;
  {SERDES, 4'd13} : slewctrl0_lane_expected = 2'b00;
  {SAS, 4'd0} : slewctrl0_lane_expected = 2'b01;
  {SAS, 4'd1} : slewctrl0_lane_expected = 2'b01;
  {SAS, 4'd2} : slewctrl0_lane_expected = 2'b01;
  {SAS, 4'd3} : slewctrl0_lane_expected = 2'b00;
  {SAS, 4'd4} : slewctrl0_lane_expected = 2'b00;
  {PCIE, 4'd0} : slewctrl0_lane_expected = 2'b01;
  {PCIE, 4'd1} : slewctrl0_lane_expected = 2'b01;
  {PCIE, 4'd2} : slewctrl0_lane_expected = 2'b00;
  {PCIE, 4'd3} : slewctrl0_lane_expected = 2'b00;
default: slewctrl0_lane_expected = 2'bzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : tx_train_pat_sel_lane_expected = 2'b00;
  {USB, 4'd2} : tx_train_pat_sel_lane_expected = 2'b00;
  {SERDES, 4'd0} : tx_train_pat_sel_lane_expected = 2'b01;
  {SERDES, 4'd1} : tx_train_pat_sel_lane_expected = 2'b01;
  {SERDES, 4'd2} : tx_train_pat_sel_lane_expected = 2'b01;
  {SERDES, 4'd3} : tx_train_pat_sel_lane_expected = 2'b01;
  {SERDES, 4'd4} : tx_train_pat_sel_lane_expected = 2'b01;
  {SERDES, 4'd5} : tx_train_pat_sel_lane_expected = 2'b01;
  {SERDES, 4'd6} : tx_train_pat_sel_lane_expected = 2'b01;
  {SERDES, 4'd7} : tx_train_pat_sel_lane_expected = 2'b10;
  {SERDES, 4'd8} : tx_train_pat_sel_lane_expected = 2'b10;
  {SERDES, 4'd9} : tx_train_pat_sel_lane_expected = 2'b10;
  {SERDES, 4'd12} : tx_train_pat_sel_lane_expected = 2'b01;
  {SERDES, 4'd13} : tx_train_pat_sel_lane_expected = 2'b10;
  {SAS, 4'd0} : tx_train_pat_sel_lane_expected = 2'b00;
  {SAS, 4'd1} : tx_train_pat_sel_lane_expected = 2'b00;
  {SAS, 4'd2} : tx_train_pat_sel_lane_expected = 2'b00;
  {SAS, 4'd3} : tx_train_pat_sel_lane_expected = 2'b00;
  {SAS, 4'd4} : tx_train_pat_sel_lane_expected = 2'b11;
  {PCIE, 4'd0} : tx_train_pat_sel_lane_expected = 2'b00;
  {PCIE, 4'd1} : tx_train_pat_sel_lane_expected = 2'b00;
  {PCIE, 4'd2} : tx_train_pat_sel_lane_expected = 2'b00;
  {PCIE, 4'd3} : tx_train_pat_sel_lane_expected = 2'b00;
default: tx_train_pat_sel_lane_expected = 2'bzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : train_pat_num_lane_expected = 9'b001000010;
  {USB, 4'd2} : train_pat_num_lane_expected = 9'b001000010;
  {SERDES, 4'd0} : train_pat_num_lane_expected = 9'b010001000;
  {SERDES, 4'd1} : train_pat_num_lane_expected = 9'b010001000;
  {SERDES, 4'd2} : train_pat_num_lane_expected = 9'b010001000;
  {SERDES, 4'd3} : train_pat_num_lane_expected = 9'b010001000;
  {SERDES, 4'd4} : train_pat_num_lane_expected = 9'b010001000;
  {SERDES, 4'd5} : train_pat_num_lane_expected = 9'b010001000;
  {SERDES, 4'd6} : train_pat_num_lane_expected = 9'b010001000;
  {SERDES, 4'd7} : train_pat_num_lane_expected = 9'b010001000;
  {SERDES, 4'd8} : train_pat_num_lane_expected = 9'b010001000;
  {SERDES, 4'd9} : train_pat_num_lane_expected = 9'b010001000;
  {SERDES, 4'd12} : train_pat_num_lane_expected = 9'b010001000;
  {SERDES, 4'd13} : train_pat_num_lane_expected = 9'b010001000;
  {SAS, 4'd0} : train_pat_num_lane_expected = 9'b001000010;
  {SAS, 4'd1} : train_pat_num_lane_expected = 9'b001000010;
  {SAS, 4'd2} : train_pat_num_lane_expected = 9'b001000010;
  {SAS, 4'd3} : train_pat_num_lane_expected = 9'b001000010;
  {SAS, 4'd4} : train_pat_num_lane_expected = 9'b011101001;
  {PCIE, 4'd0} : train_pat_num_lane_expected = 9'b001000010;
  {PCIE, 4'd1} : train_pat_num_lane_expected = 9'b001000010;
  {PCIE, 4'd2} : train_pat_num_lane_expected = 9'b001000010;
  {PCIE, 4'd3} : train_pat_num_lane_expected = 9'b001000010;
default: train_pat_num_lane_expected = 9'bzzzzzzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : tx_train_pat_toggle_lane_expected = 1'b1;
  {USB, 4'd2} : tx_train_pat_toggle_lane_expected = 1'b1;
  {SERDES, 4'd0} : tx_train_pat_toggle_lane_expected = 1'b0;
  {SERDES, 4'd1} : tx_train_pat_toggle_lane_expected = 1'b0;
  {SERDES, 4'd2} : tx_train_pat_toggle_lane_expected = 1'b0;
  {SERDES, 4'd3} : tx_train_pat_toggle_lane_expected = 1'b0;
  {SERDES, 4'd4} : tx_train_pat_toggle_lane_expected = 1'b0;
  {SERDES, 4'd5} : tx_train_pat_toggle_lane_expected = 1'b0;
  {SERDES, 4'd6} : tx_train_pat_toggle_lane_expected = 1'b0;
  {SERDES, 4'd7} : tx_train_pat_toggle_lane_expected = 1'b0;
  {SERDES, 4'd8} : tx_train_pat_toggle_lane_expected = 1'b0;
  {SERDES, 4'd9} : tx_train_pat_toggle_lane_expected = 1'b0;
  {SERDES, 4'd12} : tx_train_pat_toggle_lane_expected = 1'b0;
  {SERDES, 4'd13} : tx_train_pat_toggle_lane_expected = 1'b0;
  {SAS, 4'd0} : tx_train_pat_toggle_lane_expected = 1'b1;
  {SAS, 4'd1} : tx_train_pat_toggle_lane_expected = 1'b1;
  {SAS, 4'd2} : tx_train_pat_toggle_lane_expected = 1'b1;
  {SAS, 4'd3} : tx_train_pat_toggle_lane_expected = 1'b1;
  {SAS, 4'd4} : tx_train_pat_toggle_lane_expected = 1'b0;
  {PCIE, 4'd0} : tx_train_pat_toggle_lane_expected = 1'b1;
  {PCIE, 4'd1} : tx_train_pat_toggle_lane_expected = 1'b1;
  {PCIE, 4'd2} : tx_train_pat_toggle_lane_expected = 1'b1;
  {PCIE, 4'd3} : tx_train_pat_toggle_lane_expected = 1'b1;
default: tx_train_pat_toggle_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : packet_sync_dis_lane_expected = 1'b1;
  {USB, 4'd2} : packet_sync_dis_lane_expected = 1'b1;
  {SERDES, 4'd0} : packet_sync_dis_lane_expected = 1'b1;
  {SERDES, 4'd1} : packet_sync_dis_lane_expected = 1'b1;
  {SERDES, 4'd2} : packet_sync_dis_lane_expected = 1'b1;
  {SERDES, 4'd3} : packet_sync_dis_lane_expected = 1'b1;
  {SERDES, 4'd4} : packet_sync_dis_lane_expected = 1'b1;
  {SERDES, 4'd5} : packet_sync_dis_lane_expected = 1'b1;
  {SERDES, 4'd6} : packet_sync_dis_lane_expected = 1'b1;
  {SERDES, 4'd7} : packet_sync_dis_lane_expected = 1'b1;
  {SERDES, 4'd8} : packet_sync_dis_lane_expected = 1'b1;
  {SERDES, 4'd9} : packet_sync_dis_lane_expected = 1'b1;
  {SERDES, 4'd12} : packet_sync_dis_lane_expected = 1'b1;
  {SERDES, 4'd13} : packet_sync_dis_lane_expected = 1'b1;
  {SAS, 4'd0} : packet_sync_dis_lane_expected = 1'b1;
  {SAS, 4'd1} : packet_sync_dis_lane_expected = 1'b1;
  {SAS, 4'd2} : packet_sync_dis_lane_expected = 1'b1;
  {SAS, 4'd3} : packet_sync_dis_lane_expected = 1'b1;
  {SAS, 4'd4} : packet_sync_dis_lane_expected = 1'b0;
  {PCIE, 4'd0} : packet_sync_dis_lane_expected = 1'b1;
  {PCIE, 4'd1} : packet_sync_dis_lane_expected = 1'b1;
  {PCIE, 4'd2} : packet_sync_dis_lane_expected = 1'b1;
  {PCIE, 4'd3} : packet_sync_dis_lane_expected = 1'b1;
default: packet_sync_dis_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : sync_det_dis_lane_expected = 1'b0;
  {USB, 4'd2} : sync_det_dis_lane_expected = 1'b0;
  {SERDES, 4'd0} : sync_det_dis_lane_expected = 1'b0;
  {SERDES, 4'd1} : sync_det_dis_lane_expected = 1'b0;
  {SERDES, 4'd2} : sync_det_dis_lane_expected = 1'b0;
  {SERDES, 4'd3} : sync_det_dis_lane_expected = 1'b0;
  {SERDES, 4'd4} : sync_det_dis_lane_expected = 1'b0;
  {SERDES, 4'd5} : sync_det_dis_lane_expected = 1'b0;
  {SERDES, 4'd6} : sync_det_dis_lane_expected = 1'b0;
  {SERDES, 4'd7} : sync_det_dis_lane_expected = 1'b0;
  {SERDES, 4'd8} : sync_det_dis_lane_expected = 1'b0;
  {SERDES, 4'd9} : sync_det_dis_lane_expected = 1'b0;
  {SERDES, 4'd12} : sync_det_dis_lane_expected = 1'b0;
  {SERDES, 4'd13} : sync_det_dis_lane_expected = 1'b0;
  {SAS, 4'd0} : sync_det_dis_lane_expected = 1'b0;
  {SAS, 4'd1} : sync_det_dis_lane_expected = 1'b0;
  {SAS, 4'd2} : sync_det_dis_lane_expected = 1'b0;
  {SAS, 4'd3} : sync_det_dis_lane_expected = 1'b0;
  {SAS, 4'd4} : sync_det_dis_lane_expected = 1'b1;
  {PCIE, 4'd0} : sync_det_dis_lane_expected = 1'b0;
  {PCIE, 4'd1} : sync_det_dis_lane_expected = 1'b0;
  {PCIE, 4'd2} : sync_det_dis_lane_expected = 1'b0;
  {PCIE, 4'd3} : sync_det_dis_lane_expected = 1'b0;
default: sync_det_dis_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : pll_rate_sel_rx_expected = 4'b0000;
  {USB, 4'd2} : pll_rate_sel_rx_expected = 4'b0000;
  {SERDES, 4'd0} : pll_rate_sel_rx_expected = 4'b0000;
  {SERDES, 4'd1} : pll_rate_sel_rx_expected = 4'b0011;
  {SERDES, 4'd2} : pll_rate_sel_rx_expected = 4'b0001;
  {SERDES, 4'd3} : pll_rate_sel_rx_expected = 4'b0011;
  {SERDES, 4'd4} : pll_rate_sel_rx_expected = 4'b0001;
  {SERDES, 4'd5} : pll_rate_sel_rx_expected = 4'b0010;
  {SERDES, 4'd6} : pll_rate_sel_rx_expected = 4'b0011;
  {SERDES, 4'd7} : pll_rate_sel_rx_expected = 4'b0100;
  {SERDES, 4'd8} : pll_rate_sel_rx_expected = 4'b0101;
  {SERDES, 4'd9} : pll_rate_sel_rx_expected = 4'b0110;
  {SERDES, 4'd12} : pll_rate_sel_rx_expected = 4'b0000;
  {SERDES, 4'd13} : pll_rate_sel_rx_expected = 4'b0001;
  {SAS, 4'd0} : pll_rate_sel_rx_expected = 4'b0001;
  {SAS, 4'd1} : pll_rate_sel_rx_expected = 4'b0001;
  {SAS, 4'd2} : pll_rate_sel_rx_expected = 4'b0001;
  {SAS, 4'd3} : pll_rate_sel_rx_expected = 4'b0001;
  {SAS, 4'd4} : pll_rate_sel_rx_expected = 4'b0000;
  {PCIE, 4'd0} : pll_rate_sel_rx_expected = 4'b0001;
  {PCIE, 4'd1} : pll_rate_sel_rx_expected = 4'b0001;
  {PCIE, 4'd2} : pll_rate_sel_rx_expected = 4'b0000;
  {PCIE, 4'd3} : pll_rate_sel_rx_expected = 4'b0000;
default: pll_rate_sel_rx_expected = 4'bzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : rx_ck_sel_lane_expected = 1'b0;
  {USB, 4'd2} : rx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd0} : rx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd1} : rx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd2} : rx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd3} : rx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd4} : rx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd5} : rx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd6} : rx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd7} : rx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd8} : rx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd9} : rx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd12} : rx_ck_sel_lane_expected = 1'b0;
  {SERDES, 4'd13} : rx_ck_sel_lane_expected = 1'b0;
  {SAS, 4'd0} : rx_ck_sel_lane_expected = 1'b0;
  {SAS, 4'd1} : rx_ck_sel_lane_expected = 1'b0;
  {SAS, 4'd2} : rx_ck_sel_lane_expected = 1'b0;
  {SAS, 4'd3} : rx_ck_sel_lane_expected = 1'b0;
  {SAS, 4'd4} : rx_ck_sel_lane_expected = 1'b0;
  {PCIE, 4'd0} : rx_ck_sel_lane_expected = 1'b1;
  {PCIE, 4'd1} : rx_ck_sel_lane_expected = 1'b1;
  {PCIE, 4'd2} : rx_ck_sel_lane_expected = 1'b0;
  {PCIE, 4'd3} : rx_ck_sel_lane_expected = 1'b0;
default: rx_ck_sel_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : rx_vddcal_rate_en_lane_expected = 1'b1;
  {USB, 4'd2} : rx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd0} : rx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd1} : rx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd2} : rx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd3} : rx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd4} : rx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd5} : rx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd6} : rx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd7} : rx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd8} : rx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd9} : rx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd12} : rx_vddcal_rate_en_lane_expected = 1'b1;
  {SERDES, 4'd13} : rx_vddcal_rate_en_lane_expected = 1'b1;
  {SAS, 4'd0} : rx_vddcal_rate_en_lane_expected = 1'b1;
  {SAS, 4'd1} : rx_vddcal_rate_en_lane_expected = 1'b1;
  {SAS, 4'd2} : rx_vddcal_rate_en_lane_expected = 1'b1;
  {SAS, 4'd3} : rx_vddcal_rate_en_lane_expected = 1'b1;
  {SAS, 4'd4} : rx_vddcal_rate_en_lane_expected = 1'b1;
  {PCIE, 4'd0} : rx_vddcal_rate_en_lane_expected = 1'b1;
  {PCIE, 4'd1} : rx_vddcal_rate_en_lane_expected = 1'b1;
  {PCIE, 4'd2} : rx_vddcal_rate_en_lane_expected = 1'b1;
  {PCIE, 4'd3} : rx_vddcal_rate_en_lane_expected = 1'b1;
default: rx_vddcal_rate_en_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : rx_speed_div_lane_expected = 3'b101;
  {USB, 4'd2} : rx_speed_div_lane_expected = 3'b100;
  {SERDES, 4'd0} : rx_speed_div_lane_expected = 3'b111;
  {SERDES, 4'd1} : rx_speed_div_lane_expected = 3'b110;
  {SERDES, 4'd2} : rx_speed_div_lane_expected = 3'b101;
  {SERDES, 4'd3} : rx_speed_div_lane_expected = 3'b101;
  {SERDES, 4'd4} : rx_speed_div_lane_expected = 3'b100;
  {SERDES, 4'd5} : rx_speed_div_lane_expected = 3'b100;
  {SERDES, 4'd6} : rx_speed_div_lane_expected = 3'b100;
  {SERDES, 4'd7} : rx_speed_div_lane_expected = 3'b000;
  {SERDES, 4'd8} : rx_speed_div_lane_expected = 3'b000;
  {SERDES, 4'd9} : rx_speed_div_lane_expected = 3'b000;
  {SERDES, 4'd12} : rx_speed_div_lane_expected = 3'b110;
  {SERDES, 4'd13} : rx_speed_div_lane_expected = 3'b000;
  {SAS, 4'd0} : rx_speed_div_lane_expected = 3'b111;
  {SAS, 4'd1} : rx_speed_div_lane_expected = 3'b110;
  {SAS, 4'd2} : rx_speed_div_lane_expected = 3'b101;
  {SAS, 4'd3} : rx_speed_div_lane_expected = 3'b100;
  {SAS, 4'd4} : rx_speed_div_lane_expected = 3'b000;
  {PCIE, 4'd0} : rx_speed_div_lane_expected = 3'b110;
  {PCIE, 4'd1} : rx_speed_div_lane_expected = 3'b101;
  {PCIE, 4'd2} : rx_speed_div_lane_expected = 3'b100;
  {PCIE, 4'd3} : rx_speed_div_lane_expected = 3'b000;
default: rx_speed_div_lane_expected = 3'bzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : dtl_clk_speedup_lane_expected = 3'b001;
  {USB, 4'd2} : dtl_clk_speedup_lane_expected = 3'b000;
  {SERDES, 4'd0} : dtl_clk_speedup_lane_expected = 3'b011;
  {SERDES, 4'd1} : dtl_clk_speedup_lane_expected = 3'b010;
  {SERDES, 4'd2} : dtl_clk_speedup_lane_expected = 3'b001;
  {SERDES, 4'd3} : dtl_clk_speedup_lane_expected = 3'b001;
  {SERDES, 4'd4} : dtl_clk_speedup_lane_expected = 3'b000;
  {SERDES, 4'd5} : dtl_clk_speedup_lane_expected = 3'b000;
  {SERDES, 4'd6} : dtl_clk_speedup_lane_expected = 3'b000;
  {SERDES, 4'd7} : dtl_clk_speedup_lane_expected = 3'b100;
  {SERDES, 4'd8} : dtl_clk_speedup_lane_expected = 3'b100;
  {SERDES, 4'd9} : dtl_clk_speedup_lane_expected = 3'b100;
  {SERDES, 4'd12} : dtl_clk_speedup_lane_expected = 3'b010;
  {SERDES, 4'd13} : dtl_clk_speedup_lane_expected = 3'b100;
  {SAS, 4'd0} : dtl_clk_speedup_lane_expected = 3'b011;
  {SAS, 4'd1} : dtl_clk_speedup_lane_expected = 3'b010;
  {SAS, 4'd2} : dtl_clk_speedup_lane_expected = 3'b001;
  {SAS, 4'd3} : dtl_clk_speedup_lane_expected = 3'b000;
  {SAS, 4'd4} : dtl_clk_speedup_lane_expected = 3'b100;
  {PCIE, 4'd0} : dtl_clk_speedup_lane_expected = 3'b010;
  {PCIE, 4'd1} : dtl_clk_speedup_lane_expected = 3'b001;
  {PCIE, 4'd2} : dtl_clk_speedup_lane_expected = 3'b000;
  {PCIE, 4'd3} : dtl_clk_speedup_lane_expected = 3'b100;
default: dtl_clk_speedup_lane_expected = 3'bzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : intpi_lane_expected = 4'b1000;
  {USB, 4'd2} : intpi_lane_expected = 4'b1000;
  {SERDES, 4'd0} : intpi_lane_expected = 4'b1000;
  {SERDES, 4'd1} : intpi_lane_expected = 4'b1011;
  {SERDES, 4'd2} : intpi_lane_expected = 4'b1000;
  {SERDES, 4'd3} : intpi_lane_expected = 4'b1011;
  {SERDES, 4'd4} : intpi_lane_expected = 4'b1000;
  {SERDES, 4'd5} : intpi_lane_expected = 4'b1011;
  {SERDES, 4'd6} : intpi_lane_expected = 4'b1011;
  {SERDES, 4'd7} : intpi_lane_expected = 4'b1101;
  {SERDES, 4'd8} : intpi_lane_expected = 4'b1101;
  {SERDES, 4'd9} : intpi_lane_expected = 4'b1101;
  {SERDES, 4'd12} : intpi_lane_expected = 4'b1000;
  {SERDES, 4'd13} : intpi_lane_expected = 4'b1000;
  {SAS, 4'd0} : intpi_lane_expected = 4'b1011;
  {SAS, 4'd1} : intpi_lane_expected = 4'b1011;
  {SAS, 4'd2} : intpi_lane_expected = 4'b1011;
  {SAS, 4'd3} : intpi_lane_expected = 4'b1011;
  {SAS, 4'd4} : intpi_lane_expected = 4'b1010;
  {PCIE, 4'd0} : intpi_lane_expected = 4'b1000;
  {PCIE, 4'd1} : intpi_lane_expected = 4'b1000;
  {PCIE, 4'd2} : intpi_lane_expected = 4'b0101;
  {PCIE, 4'd3} : intpi_lane_expected = 4'b0101;
default: intpi_lane_expected = 4'bzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : intpr_lane_expected = 2'b10;
  {USB, 4'd2} : intpr_lane_expected = 2'b10;
  {SERDES, 4'd0} : intpr_lane_expected = 2'b10;
  {SERDES, 4'd1} : intpr_lane_expected = 2'b01;
  {SERDES, 4'd2} : intpr_lane_expected = 2'b10;
  {SERDES, 4'd3} : intpr_lane_expected = 2'b01;
  {SERDES, 4'd4} : intpr_lane_expected = 2'b10;
  {SERDES, 4'd5} : intpr_lane_expected = 2'b01;
  {SERDES, 4'd6} : intpr_lane_expected = 2'b01;
  {SERDES, 4'd7} : intpr_lane_expected = 2'b01;
  {SERDES, 4'd8} : intpr_lane_expected = 2'b00;
  {SERDES, 4'd9} : intpr_lane_expected = 2'b00;
  {SERDES, 4'd12} : intpr_lane_expected = 2'b10;
  {SERDES, 4'd13} : intpr_lane_expected = 2'b10;
  {SAS, 4'd0} : intpr_lane_expected = 2'b01;
  {SAS, 4'd1} : intpr_lane_expected = 2'b01;
  {SAS, 4'd2} : intpr_lane_expected = 2'b01;
  {SAS, 4'd3} : intpr_lane_expected = 2'b01;
  {SAS, 4'd4} : intpr_lane_expected = 2'b01;
  {PCIE, 4'd0} : intpr_lane_expected = 2'b10;
  {PCIE, 4'd1} : intpr_lane_expected = 2'b10;
  {PCIE, 4'd2} : intpr_lane_expected = 2'b11;
  {PCIE, 4'd3} : intpr_lane_expected = 2'b11;
default: intpr_lane_expected = 2'bzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : dll_freq_sel_lane_expected = 3'b100;
  {USB, 4'd2} : dll_freq_sel_lane_expected = 3'b100;
  {SERDES, 4'd0} : dll_freq_sel_lane_expected = 3'b100;
  {SERDES, 4'd1} : dll_freq_sel_lane_expected = 3'b110;
  {SERDES, 4'd2} : dll_freq_sel_lane_expected = 3'b100;
  {SERDES, 4'd3} : dll_freq_sel_lane_expected = 3'b110;
  {SERDES, 4'd4} : dll_freq_sel_lane_expected = 3'b100;
  {SERDES, 4'd5} : dll_freq_sel_lane_expected = 3'b110;
  {SERDES, 4'd6} : dll_freq_sel_lane_expected = 3'b110;
  {SERDES, 4'd7} : dll_freq_sel_lane_expected = 3'b110;
  {SERDES, 4'd8} : dll_freq_sel_lane_expected = 3'b110;
  {SERDES, 4'd9} : dll_freq_sel_lane_expected = 3'b110;
  {SERDES, 4'd12} : dll_freq_sel_lane_expected = 3'b100;
  {SERDES, 4'd13} : dll_freq_sel_lane_expected = 3'b100;
  {SAS, 4'd0} : dll_freq_sel_lane_expected = 3'b110;
  {SAS, 4'd1} : dll_freq_sel_lane_expected = 3'b110;
  {SAS, 4'd2} : dll_freq_sel_lane_expected = 3'b110;
  {SAS, 4'd3} : dll_freq_sel_lane_expected = 3'b110;
  {SAS, 4'd4} : dll_freq_sel_lane_expected = 3'b100;
  {PCIE, 4'd0} : dll_freq_sel_lane_expected = 3'b100;
  {PCIE, 4'd1} : dll_freq_sel_lane_expected = 3'b100;
  {PCIE, 4'd2} : dll_freq_sel_lane_expected = 3'b000;
  {PCIE, 4'd3} : dll_freq_sel_lane_expected = 3'b000;
default: dll_freq_sel_lane_expected = 3'bzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : eom_dll_freq_sel_lane_expected = 3'b100;
  {USB, 4'd2} : eom_dll_freq_sel_lane_expected = 3'b100;
  {SERDES, 4'd0} : eom_dll_freq_sel_lane_expected = 3'b100;
  {SERDES, 4'd1} : eom_dll_freq_sel_lane_expected = 3'b110;
  {SERDES, 4'd2} : eom_dll_freq_sel_lane_expected = 3'b100;
  {SERDES, 4'd3} : eom_dll_freq_sel_lane_expected = 3'b110;
  {SERDES, 4'd4} : eom_dll_freq_sel_lane_expected = 3'b100;
  {SERDES, 4'd5} : eom_dll_freq_sel_lane_expected = 3'b110;
  {SERDES, 4'd6} : eom_dll_freq_sel_lane_expected = 3'b110;
  {SERDES, 4'd7} : eom_dll_freq_sel_lane_expected = 3'b110;
  {SERDES, 4'd8} : eom_dll_freq_sel_lane_expected = 3'b110;
  {SERDES, 4'd9} : eom_dll_freq_sel_lane_expected = 3'b110;
  {SERDES, 4'd12} : eom_dll_freq_sel_lane_expected = 3'b100;
  {SERDES, 4'd13} : eom_dll_freq_sel_lane_expected = 3'b100;
  {SAS, 4'd0} : eom_dll_freq_sel_lane_expected = 3'b110;
  {SAS, 4'd1} : eom_dll_freq_sel_lane_expected = 3'b110;
  {SAS, 4'd2} : eom_dll_freq_sel_lane_expected = 3'b110;
  {SAS, 4'd3} : eom_dll_freq_sel_lane_expected = 3'b110;
  {SAS, 4'd4} : eom_dll_freq_sel_lane_expected = 3'b100;
  {PCIE, 4'd0} : eom_dll_freq_sel_lane_expected = 3'b100;
  {PCIE, 4'd1} : eom_dll_freq_sel_lane_expected = 3'b100;
  {PCIE, 4'd2} : eom_dll_freq_sel_lane_expected = 3'b000;
  {PCIE, 4'd3} : eom_dll_freq_sel_lane_expected = 3'b000;
default: eom_dll_freq_sel_lane_expected = 3'bzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : align90_8g_en_lane_expected = 1'b0;
  {USB, 4'd2} : align90_8g_en_lane_expected = 1'b0;
  {SERDES, 4'd0} : align90_8g_en_lane_expected = 1'b0;
  {SERDES, 4'd1} : align90_8g_en_lane_expected = 1'b0;
  {SERDES, 4'd2} : align90_8g_en_lane_expected = 1'b0;
  {SERDES, 4'd3} : align90_8g_en_lane_expected = 1'b0;
  {SERDES, 4'd4} : align90_8g_en_lane_expected = 1'b0;
  {SERDES, 4'd5} : align90_8g_en_lane_expected = 1'b0;
  {SERDES, 4'd6} : align90_8g_en_lane_expected = 1'b0;
  {SERDES, 4'd7} : align90_8g_en_lane_expected = 1'b0;
  {SERDES, 4'd8} : align90_8g_en_lane_expected = 1'b0;
  {SERDES, 4'd9} : align90_8g_en_lane_expected = 1'b0;
  {SERDES, 4'd12} : align90_8g_en_lane_expected = 1'b0;
  {SERDES, 4'd13} : align90_8g_en_lane_expected = 1'b0;
  {SAS, 4'd0} : align90_8g_en_lane_expected = 1'b0;
  {SAS, 4'd1} : align90_8g_en_lane_expected = 1'b0;
  {SAS, 4'd2} : align90_8g_en_lane_expected = 1'b0;
  {SAS, 4'd3} : align90_8g_en_lane_expected = 1'b0;
  {SAS, 4'd4} : align90_8g_en_lane_expected = 1'b0;
  {PCIE, 4'd0} : align90_8g_en_lane_expected = 1'b0;
  {PCIE, 4'd1} : align90_8g_en_lane_expected = 1'b0;
  {PCIE, 4'd2} : align90_8g_en_lane_expected = 1'b1;
  {PCIE, 4'd3} : align90_8g_en_lane_expected = 1'b1;
default: align90_8g_en_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : rx_reg0p9_speed_track_clk_lane_expected = 3'b001;
  {USB, 4'd2} : rx_reg0p9_speed_track_clk_lane_expected = 3'b001;
  {SERDES, 4'd0} : rx_reg0p9_speed_track_clk_lane_expected = 3'b001;
  {SERDES, 4'd1} : rx_reg0p9_speed_track_clk_lane_expected = 3'b011;
  {SERDES, 4'd2} : rx_reg0p9_speed_track_clk_lane_expected = 3'b001;
  {SERDES, 4'd3} : rx_reg0p9_speed_track_clk_lane_expected = 3'b011;
  {SERDES, 4'd4} : rx_reg0p9_speed_track_clk_lane_expected = 3'b001;
  {SERDES, 4'd5} : rx_reg0p9_speed_track_clk_lane_expected = 3'b011;
  {SERDES, 4'd6} : rx_reg0p9_speed_track_clk_lane_expected = 3'b011;
  {SERDES, 4'd7} : rx_reg0p9_speed_track_clk_lane_expected = 3'b111;
  {SERDES, 4'd8} : rx_reg0p9_speed_track_clk_lane_expected = 3'b111;
  {SERDES, 4'd9} : rx_reg0p9_speed_track_clk_lane_expected = 3'b111;
  {SERDES, 4'd12} : rx_reg0p9_speed_track_clk_lane_expected = 3'b001;
  {SERDES, 4'd13} : rx_reg0p9_speed_track_clk_lane_expected = 3'b001;
  {SAS, 4'd0} : rx_reg0p9_speed_track_clk_lane_expected = 3'b011;
  {SAS, 4'd1} : rx_reg0p9_speed_track_clk_lane_expected = 3'b011;
  {SAS, 4'd2} : rx_reg0p9_speed_track_clk_lane_expected = 3'b011;
  {SAS, 4'd3} : rx_reg0p9_speed_track_clk_lane_expected = 3'b011;
  {SAS, 4'd4} : rx_reg0p9_speed_track_clk_lane_expected = 3'b001;
  {PCIE, 4'd0} : rx_reg0p9_speed_track_clk_lane_expected = 3'b001;
  {PCIE, 4'd1} : rx_reg0p9_speed_track_clk_lane_expected = 3'b001;
  {PCIE, 4'd2} : rx_reg0p9_speed_track_clk_lane_expected = 3'b000;
  {PCIE, 4'd3} : rx_reg0p9_speed_track_clk_lane_expected = 3'b000;
default: rx_reg0p9_speed_track_clk_lane_expected = 3'bzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : rx_reg0p9_speed_track_clk_half_lane_expected = 1'b1;
  {USB, 4'd2} : rx_reg0p9_speed_track_clk_half_lane_expected = 1'b1;
  {SERDES, 4'd0} : rx_reg0p9_speed_track_clk_half_lane_expected = 1'b1;
  {SERDES, 4'd1} : rx_reg0p9_speed_track_clk_half_lane_expected = 1'b1;
  {SERDES, 4'd2} : rx_reg0p9_speed_track_clk_half_lane_expected = 1'b1;
  {SERDES, 4'd3} : rx_reg0p9_speed_track_clk_half_lane_expected = 1'b1;
  {SERDES, 4'd4} : rx_reg0p9_speed_track_clk_half_lane_expected = 1'b1;
  {SERDES, 4'd5} : rx_reg0p9_speed_track_clk_half_lane_expected = 1'b1;
  {SERDES, 4'd6} : rx_reg0p9_speed_track_clk_half_lane_expected = 1'b1;
  {SERDES, 4'd7} : rx_reg0p9_speed_track_clk_half_lane_expected = 1'b0;
  {SERDES, 4'd8} : rx_reg0p9_speed_track_clk_half_lane_expected = 1'b0;
  {SERDES, 4'd9} : rx_reg0p9_speed_track_clk_half_lane_expected = 1'b0;
  {SERDES, 4'd12} : rx_reg0p9_speed_track_clk_half_lane_expected = 1'b1;
  {SERDES, 4'd13} : rx_reg0p9_speed_track_clk_half_lane_expected = 1'b0;
  {SAS, 4'd0} : rx_reg0p9_speed_track_clk_half_lane_expected = 1'b1;
  {SAS, 4'd1} : rx_reg0p9_speed_track_clk_half_lane_expected = 1'b1;
  {SAS, 4'd2} : rx_reg0p9_speed_track_clk_half_lane_expected = 1'b1;
  {SAS, 4'd3} : rx_reg0p9_speed_track_clk_half_lane_expected = 1'b1;
  {SAS, 4'd4} : rx_reg0p9_speed_track_clk_half_lane_expected = 1'b0;
  {PCIE, 4'd0} : rx_reg0p9_speed_track_clk_half_lane_expected = 1'b1;
  {PCIE, 4'd1} : rx_reg0p9_speed_track_clk_half_lane_expected = 1'b1;
  {PCIE, 4'd2} : rx_reg0p9_speed_track_clk_half_lane_expected = 1'b1;
  {PCIE, 4'd3} : rx_reg0p9_speed_track_clk_half_lane_expected = 1'b0;
default: rx_reg0p9_speed_track_clk_half_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : rx_reg0p9_speed_track_data_lane_expected = 3'b110;
  {USB, 4'd2} : rx_reg0p9_speed_track_data_lane_expected = 3'b110;
  {SERDES, 4'd0} : rx_reg0p9_speed_track_data_lane_expected = 3'b110;
  {SERDES, 4'd1} : rx_reg0p9_speed_track_data_lane_expected = 3'b110;
  {SERDES, 4'd2} : rx_reg0p9_speed_track_data_lane_expected = 3'b110;
  {SERDES, 4'd3} : rx_reg0p9_speed_track_data_lane_expected = 3'b110;
  {SERDES, 4'd4} : rx_reg0p9_speed_track_data_lane_expected = 3'b110;
  {SERDES, 4'd5} : rx_reg0p9_speed_track_data_lane_expected = 3'b110;
  {SERDES, 4'd6} : rx_reg0p9_speed_track_data_lane_expected = 3'b110;
  {SERDES, 4'd7} : rx_reg0p9_speed_track_data_lane_expected = 3'b110;
  {SERDES, 4'd8} : rx_reg0p9_speed_track_data_lane_expected = 3'b110;
  {SERDES, 4'd9} : rx_reg0p9_speed_track_data_lane_expected = 3'b110;
  {SERDES, 4'd12} : rx_reg0p9_speed_track_data_lane_expected = 3'b110;
  {SERDES, 4'd13} : rx_reg0p9_speed_track_data_lane_expected = 3'b110;
  {SAS, 4'd0} : rx_reg0p9_speed_track_data_lane_expected = 3'b110;
  {SAS, 4'd1} : rx_reg0p9_speed_track_data_lane_expected = 3'b110;
  {SAS, 4'd2} : rx_reg0p9_speed_track_data_lane_expected = 3'b110;
  {SAS, 4'd3} : rx_reg0p9_speed_track_data_lane_expected = 3'b110;
  {SAS, 4'd4} : rx_reg0p9_speed_track_data_lane_expected = 3'b110;
  {PCIE, 4'd0} : rx_reg0p9_speed_track_data_lane_expected = 3'b110;
  {PCIE, 4'd1} : rx_reg0p9_speed_track_data_lane_expected = 3'b110;
  {PCIE, 4'd2} : rx_reg0p9_speed_track_data_lane_expected = 3'b110;
  {PCIE, 4'd3} : rx_reg0p9_speed_track_data_lane_expected = 3'b110;
default: rx_reg0p9_speed_track_data_lane_expected = 3'bzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : rx_selmufi_lane_expected = 3'b100;
  {USB, 4'd2} : rx_selmufi_lane_expected = 3'b100;
  {SERDES, 4'd0} : rx_selmufi_lane_expected = 3'b100;
  {SERDES, 4'd1} : rx_selmufi_lane_expected = 3'b100;
  {SERDES, 4'd2} : rx_selmufi_lane_expected = 3'b100;
  {SERDES, 4'd3} : rx_selmufi_lane_expected = 3'b100;
  {SERDES, 4'd4} : rx_selmufi_lane_expected = 3'b100;
  {SERDES, 4'd5} : rx_selmufi_lane_expected = 3'b100;
  {SERDES, 4'd6} : rx_selmufi_lane_expected = 3'b100;
  {SERDES, 4'd7} : rx_selmufi_lane_expected = 3'b100;
  {SERDES, 4'd8} : rx_selmufi_lane_expected = 3'b100;
  {SERDES, 4'd9} : rx_selmufi_lane_expected = 3'b100;
  {SERDES, 4'd12} : rx_selmufi_lane_expected = 3'b100;
  {SERDES, 4'd13} : rx_selmufi_lane_expected = 3'b100;
  {SAS, 4'd0} : rx_selmufi_lane_expected = 3'b100;
  {SAS, 4'd1} : rx_selmufi_lane_expected = 3'b100;
  {SAS, 4'd2} : rx_selmufi_lane_expected = 3'b100;
  {SAS, 4'd3} : rx_selmufi_lane_expected = 3'b100;
  {SAS, 4'd4} : rx_selmufi_lane_expected = 3'b100;
  {PCIE, 4'd0} : rx_selmufi_lane_expected = 3'b100;
  {PCIE, 4'd1} : rx_selmufi_lane_expected = 3'b100;
  {PCIE, 4'd2} : rx_selmufi_lane_expected = 3'b100;
  {PCIE, 4'd3} : rx_selmufi_lane_expected = 3'b100;
default: rx_selmufi_lane_expected = 3'bzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : rx_selmuff_lane_expected = 3'b100;
  {USB, 4'd2} : rx_selmuff_lane_expected = 3'b101;
  {SERDES, 4'd0} : rx_selmuff_lane_expected = 3'b101;
  {SERDES, 4'd1} : rx_selmuff_lane_expected = 3'b101;
  {SERDES, 4'd2} : rx_selmuff_lane_expected = 3'b101;
  {SERDES, 4'd3} : rx_selmuff_lane_expected = 3'b110;
  {SERDES, 4'd4} : rx_selmuff_lane_expected = 3'b101;
  {SERDES, 4'd5} : rx_selmuff_lane_expected = 3'b101;
  {SERDES, 4'd6} : rx_selmuff_lane_expected = 3'b101;
  {SERDES, 4'd7} : rx_selmuff_lane_expected = 3'b101;
  {SERDES, 4'd8} : rx_selmuff_lane_expected = 3'b101;
  {SERDES, 4'd9} : rx_selmuff_lane_expected = 3'b101;
  {SERDES, 4'd12} : rx_selmuff_lane_expected = 3'b101;
  {SERDES, 4'd13} : rx_selmuff_lane_expected = 3'b101;
  {SAS, 4'd0} : rx_selmuff_lane_expected = 3'b101;
  {SAS, 4'd1} : rx_selmuff_lane_expected = 3'b101;
  {SAS, 4'd2} : rx_selmuff_lane_expected = 3'b110;
  {SAS, 4'd3} : rx_selmuff_lane_expected = 3'b101;
  {SAS, 4'd4} : rx_selmuff_lane_expected = 3'b101;
  {PCIE, 4'd0} : rx_selmuff_lane_expected = 3'b101;
  {PCIE, 4'd1} : rx_selmuff_lane_expected = 3'b101;
  {PCIE, 4'd2} : rx_selmuff_lane_expected = 3'b101;
  {PCIE, 4'd3} : rx_selmuff_lane_expected = 3'b100;
default: rx_selmuff_lane_expected = 3'bzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : reg_selmupi_lane_expected = 4'b0011;
  {USB, 4'd2} : reg_selmupi_lane_expected = 4'b0011;
  {SERDES, 4'd0} : reg_selmupi_lane_expected = 4'b0011;
  {SERDES, 4'd1} : reg_selmupi_lane_expected = 4'b0011;
  {SERDES, 4'd2} : reg_selmupi_lane_expected = 4'b0011;
  {SERDES, 4'd3} : reg_selmupi_lane_expected = 4'b0011;
  {SERDES, 4'd4} : reg_selmupi_lane_expected = 4'b0011;
  {SERDES, 4'd5} : reg_selmupi_lane_expected = 4'b0011;
  {SERDES, 4'd6} : reg_selmupi_lane_expected = 4'b0011;
  {SERDES, 4'd7} : reg_selmupi_lane_expected = 4'b0011;
  {SERDES, 4'd8} : reg_selmupi_lane_expected = 4'b0011;
  {SERDES, 4'd9} : reg_selmupi_lane_expected = 4'b0011;
  {SERDES, 4'd12} : reg_selmupi_lane_expected = 4'b0011;
  {SERDES, 4'd13} : reg_selmupi_lane_expected = 4'b0011;
  {SAS, 4'd0} : reg_selmupi_lane_expected = 4'b0011;
  {SAS, 4'd1} : reg_selmupi_lane_expected = 4'b0011;
  {SAS, 4'd2} : reg_selmupi_lane_expected = 4'b0011;
  {SAS, 4'd3} : reg_selmupi_lane_expected = 4'b0011;
  {SAS, 4'd4} : reg_selmupi_lane_expected = 4'b0011;
  {PCIE, 4'd0} : reg_selmupi_lane_expected = 4'b0011;
  {PCIE, 4'd1} : reg_selmupi_lane_expected = 4'b0011;
  {PCIE, 4'd2} : reg_selmupi_lane_expected = 4'b0011;
  {PCIE, 4'd3} : reg_selmupi_lane_expected = 4'b0011;
default: reg_selmupi_lane_expected = 4'bzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : reg_selmupf_lane_expected = 4'b0010;
  {USB, 4'd2} : reg_selmupf_lane_expected = 4'b0100;
  {SERDES, 4'd0} : reg_selmupf_lane_expected = 4'b0010;
  {SERDES, 4'd1} : reg_selmupf_lane_expected = 4'b0010;
  {SERDES, 4'd2} : reg_selmupf_lane_expected = 4'b0010;
  {SERDES, 4'd3} : reg_selmupf_lane_expected = 4'b0010;
  {SERDES, 4'd4} : reg_selmupf_lane_expected = 4'b0100;
  {SERDES, 4'd5} : reg_selmupf_lane_expected = 4'b0011;
  {SERDES, 4'd6} : reg_selmupf_lane_expected = 4'b0011;
  {SERDES, 4'd7} : reg_selmupf_lane_expected = 4'b0100;
  {SERDES, 4'd8} : reg_selmupf_lane_expected = 4'b0100;
  {SERDES, 4'd9} : reg_selmupf_lane_expected = 4'b0100;
  {SERDES, 4'd12} : reg_selmupf_lane_expected = 4'b0010;
  {SERDES, 4'd13} : reg_selmupf_lane_expected = 4'b0100;
  {SAS, 4'd0} : reg_selmupf_lane_expected = 4'b0010;
  {SAS, 4'd1} : reg_selmupf_lane_expected = 4'b0010;
  {SAS, 4'd2} : reg_selmupf_lane_expected = 4'b0010;
  {SAS, 4'd3} : reg_selmupf_lane_expected = 4'b0011;
  {SAS, 4'd4} : reg_selmupf_lane_expected = 4'b0100;
  {PCIE, 4'd0} : reg_selmupf_lane_expected = 4'b0010;
  {PCIE, 4'd1} : reg_selmupf_lane_expected = 4'b0011;
  {PCIE, 4'd2} : reg_selmupf_lane_expected = 4'b0011;
  {PCIE, 4'd3} : reg_selmupf_lane_expected = 4'b0100;
default: reg_selmupf_lane_expected = 4'bzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : rx_rxclk_25m_ctrl_lane_expected = 2'b11;
  {USB, 4'd2} : rx_rxclk_25m_ctrl_lane_expected = 2'b11;
  {SERDES, 4'd0} : rx_rxclk_25m_ctrl_lane_expected = 2'b11;
  {SERDES, 4'd1} : rx_rxclk_25m_ctrl_lane_expected = 2'b01;
  {SERDES, 4'd2} : rx_rxclk_25m_ctrl_lane_expected = 2'b01;
  {SERDES, 4'd3} : rx_rxclk_25m_ctrl_lane_expected = 2'b01;
  {SERDES, 4'd4} : rx_rxclk_25m_ctrl_lane_expected = 2'b01;
  {SERDES, 4'd5} : rx_rxclk_25m_ctrl_lane_expected = 2'b01;
  {SERDES, 4'd6} : rx_rxclk_25m_ctrl_lane_expected = 2'b01;
  {SERDES, 4'd7} : rx_rxclk_25m_ctrl_lane_expected = 2'b11;
  {SERDES, 4'd8} : rx_rxclk_25m_ctrl_lane_expected = 2'b01;
  {SERDES, 4'd9} : rx_rxclk_25m_ctrl_lane_expected = 2'b01;
  {SERDES, 4'd12} : rx_rxclk_25m_ctrl_lane_expected = 2'b11;
  {SERDES, 4'd13} : rx_rxclk_25m_ctrl_lane_expected = 2'b01;
  {SAS, 4'd0} : rx_rxclk_25m_ctrl_lane_expected = 2'b11;
  {SAS, 4'd1} : rx_rxclk_25m_ctrl_lane_expected = 2'b11;
  {SAS, 4'd2} : rx_rxclk_25m_ctrl_lane_expected = 2'b11;
  {SAS, 4'd3} : rx_rxclk_25m_ctrl_lane_expected = 2'b11;
  {SAS, 4'd4} : rx_rxclk_25m_ctrl_lane_expected = 2'b11;
  {PCIE, 4'd0} : rx_rxclk_25m_ctrl_lane_expected = 2'b11;
  {PCIE, 4'd1} : rx_rxclk_25m_ctrl_lane_expected = 2'b11;
  {PCIE, 4'd2} : rx_rxclk_25m_ctrl_lane_expected = 2'b11;
  {PCIE, 4'd3} : rx_rxclk_25m_ctrl_lane_expected = 2'b11;
default: rx_rxclk_25m_ctrl_lane_expected = 2'bzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : rx_rxclk_25m_div1p5_en_lane_expected = 1'b0;
  {USB, 4'd2} : rx_rxclk_25m_div1p5_en_lane_expected = 1'b0;
  {SERDES, 4'd0} : rx_rxclk_25m_div1p5_en_lane_expected = 1'b0;
  {SERDES, 4'd1} : rx_rxclk_25m_div1p5_en_lane_expected = 1'b0;
  {SERDES, 4'd2} : rx_rxclk_25m_div1p5_en_lane_expected = 1'b1;
  {SERDES, 4'd3} : rx_rxclk_25m_div1p5_en_lane_expected = 1'b0;
  {SERDES, 4'd4} : rx_rxclk_25m_div1p5_en_lane_expected = 1'b1;
  {SERDES, 4'd5} : rx_rxclk_25m_div1p5_en_lane_expected = 1'b1;
  {SERDES, 4'd6} : rx_rxclk_25m_div1p5_en_lane_expected = 1'b0;
  {SERDES, 4'd7} : rx_rxclk_25m_div1p5_en_lane_expected = 1'b1;
  {SERDES, 4'd8} : rx_rxclk_25m_div1p5_en_lane_expected = 1'b0;
  {SERDES, 4'd9} : rx_rxclk_25m_div1p5_en_lane_expected = 1'b1;
  {SERDES, 4'd12} : rx_rxclk_25m_div1p5_en_lane_expected = 1'b0;
  {SERDES, 4'd13} : rx_rxclk_25m_div1p5_en_lane_expected = 1'b1;
  {SAS, 4'd0} : rx_rxclk_25m_div1p5_en_lane_expected = 1'b0;
  {SAS, 4'd1} : rx_rxclk_25m_div1p5_en_lane_expected = 1'b0;
  {SAS, 4'd2} : rx_rxclk_25m_div1p5_en_lane_expected = 1'b0;
  {SAS, 4'd3} : rx_rxclk_25m_div1p5_en_lane_expected = 1'b0;
  {SAS, 4'd4} : rx_rxclk_25m_div1p5_en_lane_expected = 1'b1;
  {PCIE, 4'd0} : rx_rxclk_25m_div1p5_en_lane_expected = 1'b0;
  {PCIE, 4'd1} : rx_rxclk_25m_div1p5_en_lane_expected = 1'b0;
  {PCIE, 4'd2} : rx_rxclk_25m_div1p5_en_lane_expected = 1'b0;
  {PCIE, 4'd3} : rx_rxclk_25m_div1p5_en_lane_expected = 1'b0;
default: rx_rxclk_25m_div1p5_en_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : rx_rxclk_25m_div_lane_expected = 8'b00110010;
  {USB, 4'd2} : rx_rxclk_25m_div_lane_expected = 8'b00110010;
  {SERDES, 4'd0} : rx_rxclk_25m_div_lane_expected = 8'b00110010;
  {SERDES, 4'd1} : rx_rxclk_25m_div_lane_expected = 8'b01111101;
  {SERDES, 4'd2} : rx_rxclk_25m_div_lane_expected = 8'b10001001;
  {SERDES, 4'd3} : rx_rxclk_25m_div_lane_expected = 8'b01111101;
  {SERDES, 4'd4} : rx_rxclk_25m_div_lane_expected = 8'b10001001;
  {SERDES, 4'd5} : rx_rxclk_25m_div_lane_expected = 8'b10100010;
  {SERDES, 4'd6} : rx_rxclk_25m_div_lane_expected = 8'b01111101;
  {SERDES, 4'd7} : rx_rxclk_25m_div_lane_expected = 8'b01010110;
  {SERDES, 4'd8} : rx_rxclk_25m_div_lane_expected = 8'b10001001;
  {SERDES, 4'd9} : rx_rxclk_25m_div_lane_expected = 8'b10111011;
  {SERDES, 4'd12} : rx_rxclk_25m_div_lane_expected = 8'b00110010;
  {SERDES, 4'd13} : rx_rxclk_25m_div_lane_expected = 8'b10001001;
  {SAS, 4'd0} : rx_rxclk_25m_div_lane_expected = 8'b00111100;
  {SAS, 4'd1} : rx_rxclk_25m_div_lane_expected = 8'b00111100;
  {SAS, 4'd2} : rx_rxclk_25m_div_lane_expected = 8'b00111100;
  {SAS, 4'd3} : rx_rxclk_25m_div_lane_expected = 8'b00111100;
  {SAS, 4'd4} : rx_rxclk_25m_div_lane_expected = 8'b01001011;
  {PCIE, 4'd0} : rx_rxclk_25m_div_lane_expected = 8'b00110010;
  {PCIE, 4'd1} : rx_rxclk_25m_div_lane_expected = 8'b00110010;
  {PCIE, 4'd2} : rx_rxclk_25m_div_lane_expected = 8'b00101000;
  {PCIE, 4'd3} : rx_rxclk_25m_div_lane_expected = 8'b00101000;
default: rx_rxclk_25m_div_lane_expected = 8'bzzzzzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : rx_rxclk_25m_fix_div_en_lane_expected = 1'b1;
  {USB, 4'd2} : rx_rxclk_25m_fix_div_en_lane_expected = 1'b1;
  {SERDES, 4'd0} : rx_rxclk_25m_fix_div_en_lane_expected = 1'b1;
  {SERDES, 4'd1} : rx_rxclk_25m_fix_div_en_lane_expected = 1'b1;
  {SERDES, 4'd2} : rx_rxclk_25m_fix_div_en_lane_expected = 1'b0;
  {SERDES, 4'd3} : rx_rxclk_25m_fix_div_en_lane_expected = 1'b1;
  {SERDES, 4'd4} : rx_rxclk_25m_fix_div_en_lane_expected = 1'b0;
  {SERDES, 4'd5} : rx_rxclk_25m_fix_div_en_lane_expected = 1'b0;
  {SERDES, 4'd6} : rx_rxclk_25m_fix_div_en_lane_expected = 1'b1;
  {SERDES, 4'd7} : rx_rxclk_25m_fix_div_en_lane_expected = 1'b1;
  {SERDES, 4'd8} : rx_rxclk_25m_fix_div_en_lane_expected = 1'b0;
  {SERDES, 4'd9} : rx_rxclk_25m_fix_div_en_lane_expected = 1'b0;
  {SERDES, 4'd12} : rx_rxclk_25m_fix_div_en_lane_expected = 1'b1;
  {SERDES, 4'd13} : rx_rxclk_25m_fix_div_en_lane_expected = 1'b0;
  {SAS, 4'd0} : rx_rxclk_25m_fix_div_en_lane_expected = 1'b1;
  {SAS, 4'd1} : rx_rxclk_25m_fix_div_en_lane_expected = 1'b1;
  {SAS, 4'd2} : rx_rxclk_25m_fix_div_en_lane_expected = 1'b1;
  {SAS, 4'd3} : rx_rxclk_25m_fix_div_en_lane_expected = 1'b1;
  {SAS, 4'd4} : rx_rxclk_25m_fix_div_en_lane_expected = 1'b1;
  {PCIE, 4'd0} : rx_rxclk_25m_fix_div_en_lane_expected = 1'b1;
  {PCIE, 4'd1} : rx_rxclk_25m_fix_div_en_lane_expected = 1'b1;
  {PCIE, 4'd2} : rx_rxclk_25m_fix_div_en_lane_expected = 1'b1;
  {PCIE, 4'd3} : rx_rxclk_25m_fix_div_en_lane_expected = 1'b1;
default: rx_rxclk_25m_fix_div_en_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : dtl_clk_mode_lane_expected = 2'b10;
  {USB, 4'd2} : dtl_clk_mode_lane_expected = 2'b10;
  {SERDES, 4'd0} : dtl_clk_mode_lane_expected = 2'b10;
  {SERDES, 4'd1} : dtl_clk_mode_lane_expected = 2'b10;
  {SERDES, 4'd2} : dtl_clk_mode_lane_expected = 2'b10;
  {SERDES, 4'd3} : dtl_clk_mode_lane_expected = 2'b10;
  {SERDES, 4'd4} : dtl_clk_mode_lane_expected = 2'b10;
  {SERDES, 4'd5} : dtl_clk_mode_lane_expected = 2'b10;
  {SERDES, 4'd6} : dtl_clk_mode_lane_expected = 2'b10;
  {SERDES, 4'd7} : dtl_clk_mode_lane_expected = 2'b10;
  {SERDES, 4'd8} : dtl_clk_mode_lane_expected = 2'b10;
  {SERDES, 4'd9} : dtl_clk_mode_lane_expected = 2'b10;
  {SERDES, 4'd12} : dtl_clk_mode_lane_expected = 2'b10;
  {SERDES, 4'd13} : dtl_clk_mode_lane_expected = 2'b10;
  {SAS, 4'd0} : dtl_clk_mode_lane_expected = 2'b10;
  {SAS, 4'd1} : dtl_clk_mode_lane_expected = 2'b10;
  {SAS, 4'd2} : dtl_clk_mode_lane_expected = 2'b10;
  {SAS, 4'd3} : dtl_clk_mode_lane_expected = 2'b10;
  {SAS, 4'd4} : dtl_clk_mode_lane_expected = 2'b10;
  {PCIE, 4'd0} : dtl_clk_mode_lane_expected = 2'b10;
  {PCIE, 4'd1} : dtl_clk_mode_lane_expected = 2'b10;
  {PCIE, 4'd2} : dtl_clk_mode_lane_expected = 2'b10;
  {PCIE, 4'd3} : dtl_clk_mode_lane_expected = 2'b10;
default: dtl_clk_mode_lane_expected = 2'bzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : rx_foffset_extra_m_lane_expected = 14'b01010100001010;
  {USB, 4'd2} : rx_foffset_extra_m_lane_expected = 14'b01010100001010;
  {SERDES, 4'd0} : rx_foffset_extra_m_lane_expected = 14'b01010100001010;
  {SERDES, 4'd1} : rx_foffset_extra_m_lane_expected = 14'b01101001001101;
  {SERDES, 4'd2} : rx_foffset_extra_m_lane_expected = 14'b01010110110011;
  {SERDES, 4'd3} : rx_foffset_extra_m_lane_expected = 14'b01101001001101;
  {SERDES, 4'd4} : rx_foffset_extra_m_lane_expected = 14'b01010110110011;
  {SERDES, 4'd5} : rx_foffset_extra_m_lane_expected = 14'b01100110100101;
  {SERDES, 4'd6} : rx_foffset_extra_m_lane_expected = 14'b01101001001101;
  {SERDES, 4'd7} : rx_foffset_extra_m_lane_expected = 14'b01101100100000;
  {SERDES, 4'd8} : rx_foffset_extra_m_lane_expected = 14'b01110011101111;
  {SERDES, 4'd9} : rx_foffset_extra_m_lane_expected = 14'b01110110010111;
  {SERDES, 4'd12} : rx_foffset_extra_m_lane_expected = 14'b01010100001010;
  {SERDES, 4'd13} : rx_foffset_extra_m_lane_expected = 14'b01010110110011;
  {SAS, 4'd0} : rx_foffset_extra_m_lane_expected = 14'b01100101000000;
  {SAS, 4'd1} : rx_foffset_extra_m_lane_expected = 14'b01100101000000;
  {SAS, 4'd2} : rx_foffset_extra_m_lane_expected = 14'b01100101000000;
  {SAS, 4'd3} : rx_foffset_extra_m_lane_expected = 14'b01100101000000;
  {SAS, 4'd4} : rx_foffset_extra_m_lane_expected = 14'b01011110101100;
  {PCIE, 4'd0} : rx_foffset_extra_m_lane_expected = 14'b01010100001010;
  {PCIE, 4'd1} : rx_foffset_extra_m_lane_expected = 14'b01010100001010;
  {PCIE, 4'd2} : rx_foffset_extra_m_lane_expected = 14'b01000011010101;
  {PCIE, 4'd3} : rx_foffset_extra_m_lane_expected = 14'b01000011010101;
default: rx_foffset_extra_m_lane_expected = 14'bzzzzzzzzzzzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : init_rxfoffs_lane_expected = 10'b0000000000;
  {USB, 4'd2} : init_rxfoffs_lane_expected = 10'b0000000000;
  {SERDES, 4'd0} : init_rxfoffs_lane_expected = 10'b0000000000;
  {SERDES, 4'd1} : init_rxfoffs_lane_expected = 10'b0000000000;
  {SERDES, 4'd2} : init_rxfoffs_lane_expected = 10'b0000000000;
  {SERDES, 4'd3} : init_rxfoffs_lane_expected = 10'b0000000000;
  {SERDES, 4'd4} : init_rxfoffs_lane_expected = 10'b0000000000;
  {SERDES, 4'd5} : init_rxfoffs_lane_expected = 10'b0000000000;
  {SERDES, 4'd6} : init_rxfoffs_lane_expected = 10'b0000000000;
  {SERDES, 4'd7} : init_rxfoffs_lane_expected = 10'b0000000000;
  {SERDES, 4'd8} : init_rxfoffs_lane_expected = 10'b0000000000;
  {SERDES, 4'd9} : init_rxfoffs_lane_expected = 10'b0000000000;
  {SERDES, 4'd12} : init_rxfoffs_lane_expected = 10'b0000000000;
  {SERDES, 4'd13} : init_rxfoffs_lane_expected = 10'b0000000000;
  {SAS, 4'd0} : init_rxfoffs_lane_expected = 10'b0000000000;
  {SAS, 4'd1} : init_rxfoffs_lane_expected = 10'b0000000000;
  {SAS, 4'd2} : init_rxfoffs_lane_expected = 10'b0000000000;
  {SAS, 4'd3} : init_rxfoffs_lane_expected = 10'b0000000000;
  {SAS, 4'd4} : init_rxfoffs_lane_expected = 10'b0000000000;
  {PCIE, 4'd0} : init_rxfoffs_lane_expected = 10'b0000000000;
  {PCIE, 4'd1} : init_rxfoffs_lane_expected = 10'b0000000000;
  {PCIE, 4'd2} : init_rxfoffs_lane_expected = 10'b0000000000;
  {PCIE, 4'd3} : init_rxfoffs_lane_expected = 10'b0000000000;
default: init_rxfoffs_lane_expected = 10'bzzzzzzzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : pu_f1p_d_e_lane_expected = 1'b1;
  {USB, 4'd2} : pu_f1p_d_e_lane_expected = 1'b1;
  {SERDES, 4'd0} : pu_f1p_d_e_lane_expected = 1'b0;
  {SERDES, 4'd1} : pu_f1p_d_e_lane_expected = 1'b1;
  {SERDES, 4'd2} : pu_f1p_d_e_lane_expected = 1'b1;
  {SERDES, 4'd3} : pu_f1p_d_e_lane_expected = 1'b1;
  {SERDES, 4'd4} : pu_f1p_d_e_lane_expected = 1'b1;
  {SERDES, 4'd5} : pu_f1p_d_e_lane_expected = 1'b1;
  {SERDES, 4'd6} : pu_f1p_d_e_lane_expected = 1'b1;
  {SERDES, 4'd7} : pu_f1p_d_e_lane_expected = 1'b1;
  {SERDES, 4'd8} : pu_f1p_d_e_lane_expected = 1'b1;
  {SERDES, 4'd9} : pu_f1p_d_e_lane_expected = 1'b1;
  {SERDES, 4'd12} : pu_f1p_d_e_lane_expected = 1'b1;
  {SERDES, 4'd13} : pu_f1p_d_e_lane_expected = 1'b1;
  {SAS, 4'd0} : pu_f1p_d_e_lane_expected = 1'b0;
  {SAS, 4'd1} : pu_f1p_d_e_lane_expected = 1'b1;
  {SAS, 4'd2} : pu_f1p_d_e_lane_expected = 1'b1;
  {SAS, 4'd3} : pu_f1p_d_e_lane_expected = 1'b1;
  {SAS, 4'd4} : pu_f1p_d_e_lane_expected = 1'b1;
  {PCIE, 4'd0} : pu_f1p_d_e_lane_expected = 1'b1;
  {PCIE, 4'd1} : pu_f1p_d_e_lane_expected = 1'b1;
  {PCIE, 4'd2} : pu_f1p_d_e_lane_expected = 1'b1;
  {PCIE, 4'd3} : pu_f1p_d_e_lane_expected = 1'b1;
default: pu_f1p_d_e_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : pu_f1n_d_e_lane_expected = 1'b0;
  {USB, 4'd2} : pu_f1n_d_e_lane_expected = 1'b1;
  {SERDES, 4'd0} : pu_f1n_d_e_lane_expected = 1'b0;
  {SERDES, 4'd1} : pu_f1n_d_e_lane_expected = 1'b0;
  {SERDES, 4'd2} : pu_f1n_d_e_lane_expected = 1'b0;
  {SERDES, 4'd3} : pu_f1n_d_e_lane_expected = 1'b0;
  {SERDES, 4'd4} : pu_f1n_d_e_lane_expected = 1'b1;
  {SERDES, 4'd5} : pu_f1n_d_e_lane_expected = 1'b1;
  {SERDES, 4'd6} : pu_f1n_d_e_lane_expected = 1'b1;
  {SERDES, 4'd7} : pu_f1n_d_e_lane_expected = 1'b1;
  {SERDES, 4'd8} : pu_f1n_d_e_lane_expected = 1'b1;
  {SERDES, 4'd9} : pu_f1n_d_e_lane_expected = 1'b1;
  {SERDES, 4'd12} : pu_f1n_d_e_lane_expected = 1'b0;
  {SERDES, 4'd13} : pu_f1n_d_e_lane_expected = 1'b1;
  {SAS, 4'd0} : pu_f1n_d_e_lane_expected = 1'b0;
  {SAS, 4'd1} : pu_f1n_d_e_lane_expected = 1'b0;
  {SAS, 4'd2} : pu_f1n_d_e_lane_expected = 1'b0;
  {SAS, 4'd3} : pu_f1n_d_e_lane_expected = 1'b1;
  {SAS, 4'd4} : pu_f1n_d_e_lane_expected = 1'b1;
  {PCIE, 4'd0} : pu_f1n_d_e_lane_expected = 1'b0;
  {PCIE, 4'd1} : pu_f1n_d_e_lane_expected = 1'b0;
  {PCIE, 4'd2} : pu_f1n_d_e_lane_expected = 1'b1;
  {PCIE, 4'd3} : pu_f1n_d_e_lane_expected = 1'b1;
default: pu_f1n_d_e_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : pu_f1p_s_e_lane_expected = 1'b0;
  {USB, 4'd2} : pu_f1p_s_e_lane_expected = 1'b1;
  {SERDES, 4'd0} : pu_f1p_s_e_lane_expected = 1'b0;
  {SERDES, 4'd1} : pu_f1p_s_e_lane_expected = 1'b0;
  {SERDES, 4'd2} : pu_f1p_s_e_lane_expected = 1'b0;
  {SERDES, 4'd3} : pu_f1p_s_e_lane_expected = 1'b0;
  {SERDES, 4'd4} : pu_f1p_s_e_lane_expected = 1'b1;
  {SERDES, 4'd5} : pu_f1p_s_e_lane_expected = 1'b1;
  {SERDES, 4'd6} : pu_f1p_s_e_lane_expected = 1'b1;
  {SERDES, 4'd7} : pu_f1p_s_e_lane_expected = 1'b1;
  {SERDES, 4'd8} : pu_f1p_s_e_lane_expected = 1'b1;
  {SERDES, 4'd9} : pu_f1p_s_e_lane_expected = 1'b1;
  {SERDES, 4'd12} : pu_f1p_s_e_lane_expected = 1'b0;
  {SERDES, 4'd13} : pu_f1p_s_e_lane_expected = 1'b1;
  {SAS, 4'd0} : pu_f1p_s_e_lane_expected = 1'b0;
  {SAS, 4'd1} : pu_f1p_s_e_lane_expected = 1'b0;
  {SAS, 4'd2} : pu_f1p_s_e_lane_expected = 1'b0;
  {SAS, 4'd3} : pu_f1p_s_e_lane_expected = 1'b1;
  {SAS, 4'd4} : pu_f1p_s_e_lane_expected = 1'b1;
  {PCIE, 4'd0} : pu_f1p_s_e_lane_expected = 1'b0;
  {PCIE, 4'd1} : pu_f1p_s_e_lane_expected = 1'b0;
  {PCIE, 4'd2} : pu_f1p_s_e_lane_expected = 1'b1;
  {PCIE, 4'd3} : pu_f1p_s_e_lane_expected = 1'b1;
default: pu_f1p_s_e_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : pu_f1n_s_e_lane_expected = 1'b0;
  {USB, 4'd2} : pu_f1n_s_e_lane_expected = 1'b1;
  {SERDES, 4'd0} : pu_f1n_s_e_lane_expected = 1'b0;
  {SERDES, 4'd1} : pu_f1n_s_e_lane_expected = 1'b0;
  {SERDES, 4'd2} : pu_f1n_s_e_lane_expected = 1'b0;
  {SERDES, 4'd3} : pu_f1n_s_e_lane_expected = 1'b0;
  {SERDES, 4'd4} : pu_f1n_s_e_lane_expected = 1'b1;
  {SERDES, 4'd5} : pu_f1n_s_e_lane_expected = 1'b1;
  {SERDES, 4'd6} : pu_f1n_s_e_lane_expected = 1'b1;
  {SERDES, 4'd7} : pu_f1n_s_e_lane_expected = 1'b1;
  {SERDES, 4'd8} : pu_f1n_s_e_lane_expected = 1'b1;
  {SERDES, 4'd9} : pu_f1n_s_e_lane_expected = 1'b1;
  {SERDES, 4'd12} : pu_f1n_s_e_lane_expected = 1'b0;
  {SERDES, 4'd13} : pu_f1n_s_e_lane_expected = 1'b1;
  {SAS, 4'd0} : pu_f1n_s_e_lane_expected = 1'b0;
  {SAS, 4'd1} : pu_f1n_s_e_lane_expected = 1'b0;
  {SAS, 4'd2} : pu_f1n_s_e_lane_expected = 1'b0;
  {SAS, 4'd3} : pu_f1n_s_e_lane_expected = 1'b1;
  {SAS, 4'd4} : pu_f1n_s_e_lane_expected = 1'b1;
  {PCIE, 4'd0} : pu_f1n_s_e_lane_expected = 1'b0;
  {PCIE, 4'd1} : pu_f1n_s_e_lane_expected = 1'b0;
  {PCIE, 4'd2} : pu_f1n_s_e_lane_expected = 1'b1;
  {PCIE, 4'd3} : pu_f1n_s_e_lane_expected = 1'b1;
default: pu_f1n_s_e_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : pu_f1p_d_o_lane_expected = 1'b1;
  {USB, 4'd2} : pu_f1p_d_o_lane_expected = 1'b1;
  {SERDES, 4'd0} : pu_f1p_d_o_lane_expected = 1'b1;
  {SERDES, 4'd1} : pu_f1p_d_o_lane_expected = 1'b0;
  {SERDES, 4'd2} : pu_f1p_d_o_lane_expected = 1'b1;
  {SERDES, 4'd3} : pu_f1p_d_o_lane_expected = 1'b1;
  {SERDES, 4'd4} : pu_f1p_d_o_lane_expected = 1'b1;
  {SERDES, 4'd5} : pu_f1p_d_o_lane_expected = 1'b1;
  {SERDES, 4'd6} : pu_f1p_d_o_lane_expected = 1'b1;
  {SERDES, 4'd7} : pu_f1p_d_o_lane_expected = 1'b1;
  {SERDES, 4'd8} : pu_f1p_d_o_lane_expected = 1'b1;
  {SERDES, 4'd9} : pu_f1p_d_o_lane_expected = 1'b1;
  {SERDES, 4'd12} : pu_f1p_d_o_lane_expected = 1'b0;
  {SERDES, 4'd13} : pu_f1p_d_o_lane_expected = 1'b1;
  {SAS, 4'd0} : pu_f1p_d_o_lane_expected = 1'b1;
  {SAS, 4'd1} : pu_f1p_d_o_lane_expected = 1'b0;
  {SAS, 4'd2} : pu_f1p_d_o_lane_expected = 1'b1;
  {SAS, 4'd3} : pu_f1p_d_o_lane_expected = 1'b1;
  {SAS, 4'd4} : pu_f1p_d_o_lane_expected = 1'b1;
  {PCIE, 4'd0} : pu_f1p_d_o_lane_expected = 1'b0;
  {PCIE, 4'd1} : pu_f1p_d_o_lane_expected = 1'b1;
  {PCIE, 4'd2} : pu_f1p_d_o_lane_expected = 1'b1;
  {PCIE, 4'd3} : pu_f1p_d_o_lane_expected = 1'b1;
default: pu_f1p_d_o_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : pu_f1n_d_o_lane_expected = 1'b0;
  {USB, 4'd2} : pu_f1n_d_o_lane_expected = 1'b1;
  {SERDES, 4'd0} : pu_f1n_d_o_lane_expected = 1'b0;
  {SERDES, 4'd1} : pu_f1n_d_o_lane_expected = 1'b0;
  {SERDES, 4'd2} : pu_f1n_d_o_lane_expected = 1'b0;
  {SERDES, 4'd3} : pu_f1n_d_o_lane_expected = 1'b0;
  {SERDES, 4'd4} : pu_f1n_d_o_lane_expected = 1'b1;
  {SERDES, 4'd5} : pu_f1n_d_o_lane_expected = 1'b1;
  {SERDES, 4'd6} : pu_f1n_d_o_lane_expected = 1'b1;
  {SERDES, 4'd7} : pu_f1n_d_o_lane_expected = 1'b1;
  {SERDES, 4'd8} : pu_f1n_d_o_lane_expected = 1'b1;
  {SERDES, 4'd9} : pu_f1n_d_o_lane_expected = 1'b1;
  {SERDES, 4'd12} : pu_f1n_d_o_lane_expected = 1'b0;
  {SERDES, 4'd13} : pu_f1n_d_o_lane_expected = 1'b1;
  {SAS, 4'd0} : pu_f1n_d_o_lane_expected = 1'b0;
  {SAS, 4'd1} : pu_f1n_d_o_lane_expected = 1'b0;
  {SAS, 4'd2} : pu_f1n_d_o_lane_expected = 1'b0;
  {SAS, 4'd3} : pu_f1n_d_o_lane_expected = 1'b1;
  {SAS, 4'd4} : pu_f1n_d_o_lane_expected = 1'b1;
  {PCIE, 4'd0} : pu_f1n_d_o_lane_expected = 1'b0;
  {PCIE, 4'd1} : pu_f1n_d_o_lane_expected = 1'b0;
  {PCIE, 4'd2} : pu_f1n_d_o_lane_expected = 1'b1;
  {PCIE, 4'd3} : pu_f1n_d_o_lane_expected = 1'b1;
default: pu_f1n_d_o_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : pu_f1p_s_o_lane_expected = 1'b1;
  {USB, 4'd2} : pu_f1p_s_o_lane_expected = 1'b1;
  {SERDES, 4'd0} : pu_f1p_s_o_lane_expected = 1'b0;
  {SERDES, 4'd1} : pu_f1p_s_o_lane_expected = 1'b0;
  {SERDES, 4'd2} : pu_f1p_s_o_lane_expected = 1'b1;
  {SERDES, 4'd3} : pu_f1p_s_o_lane_expected = 1'b1;
  {SERDES, 4'd4} : pu_f1p_s_o_lane_expected = 1'b1;
  {SERDES, 4'd5} : pu_f1p_s_o_lane_expected = 1'b1;
  {SERDES, 4'd6} : pu_f1p_s_o_lane_expected = 1'b1;
  {SERDES, 4'd7} : pu_f1p_s_o_lane_expected = 1'b1;
  {SERDES, 4'd8} : pu_f1p_s_o_lane_expected = 1'b1;
  {SERDES, 4'd9} : pu_f1p_s_o_lane_expected = 1'b1;
  {SERDES, 4'd12} : pu_f1p_s_o_lane_expected = 1'b0;
  {SERDES, 4'd13} : pu_f1p_s_o_lane_expected = 1'b1;
  {SAS, 4'd0} : pu_f1p_s_o_lane_expected = 1'b0;
  {SAS, 4'd1} : pu_f1p_s_o_lane_expected = 1'b0;
  {SAS, 4'd2} : pu_f1p_s_o_lane_expected = 1'b1;
  {SAS, 4'd3} : pu_f1p_s_o_lane_expected = 1'b1;
  {SAS, 4'd4} : pu_f1p_s_o_lane_expected = 1'b1;
  {PCIE, 4'd0} : pu_f1p_s_o_lane_expected = 1'b0;
  {PCIE, 4'd1} : pu_f1p_s_o_lane_expected = 1'b1;
  {PCIE, 4'd2} : pu_f1p_s_o_lane_expected = 1'b1;
  {PCIE, 4'd3} : pu_f1p_s_o_lane_expected = 1'b1;
default: pu_f1p_s_o_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : pu_f1n_s_o_lane_expected = 1'b0;
  {USB, 4'd2} : pu_f1n_s_o_lane_expected = 1'b1;
  {SERDES, 4'd0} : pu_f1n_s_o_lane_expected = 1'b0;
  {SERDES, 4'd1} : pu_f1n_s_o_lane_expected = 1'b0;
  {SERDES, 4'd2} : pu_f1n_s_o_lane_expected = 1'b0;
  {SERDES, 4'd3} : pu_f1n_s_o_lane_expected = 1'b0;
  {SERDES, 4'd4} : pu_f1n_s_o_lane_expected = 1'b1;
  {SERDES, 4'd5} : pu_f1n_s_o_lane_expected = 1'b1;
  {SERDES, 4'd6} : pu_f1n_s_o_lane_expected = 1'b1;
  {SERDES, 4'd7} : pu_f1n_s_o_lane_expected = 1'b1;
  {SERDES, 4'd8} : pu_f1n_s_o_lane_expected = 1'b1;
  {SERDES, 4'd9} : pu_f1n_s_o_lane_expected = 1'b1;
  {SERDES, 4'd12} : pu_f1n_s_o_lane_expected = 1'b0;
  {SERDES, 4'd13} : pu_f1n_s_o_lane_expected = 1'b1;
  {SAS, 4'd0} : pu_f1n_s_o_lane_expected = 1'b0;
  {SAS, 4'd1} : pu_f1n_s_o_lane_expected = 1'b0;
  {SAS, 4'd2} : pu_f1n_s_o_lane_expected = 1'b0;
  {SAS, 4'd3} : pu_f1n_s_o_lane_expected = 1'b1;
  {SAS, 4'd4} : pu_f1n_s_o_lane_expected = 1'b1;
  {PCIE, 4'd0} : pu_f1n_s_o_lane_expected = 1'b0;
  {PCIE, 4'd1} : pu_f1n_s_o_lane_expected = 1'b0;
  {PCIE, 4'd2} : pu_f1n_s_o_lane_expected = 1'b1;
  {PCIE, 4'd3} : pu_f1n_s_o_lane_expected = 1'b1;
default: pu_f1n_s_o_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : path_disable_edge_lane_expected = 1'b1;
  {USB, 4'd2} : path_disable_edge_lane_expected = 1'b0;
  {SERDES, 4'd0} : path_disable_edge_lane_expected = 1'b1;
  {SERDES, 4'd1} : path_disable_edge_lane_expected = 1'b1;
  {SERDES, 4'd2} : path_disable_edge_lane_expected = 1'b1;
  {SERDES, 4'd3} : path_disable_edge_lane_expected = 1'b1;
  {SERDES, 4'd4} : path_disable_edge_lane_expected = 1'b0;
  {SERDES, 4'd5} : path_disable_edge_lane_expected = 1'b0;
  {SERDES, 4'd6} : path_disable_edge_lane_expected = 1'b0;
  {SERDES, 4'd7} : path_disable_edge_lane_expected = 1'b0;
  {SERDES, 4'd8} : path_disable_edge_lane_expected = 1'b0;
  {SERDES, 4'd9} : path_disable_edge_lane_expected = 1'b0;
  {SERDES, 4'd12} : path_disable_edge_lane_expected = 1'b1;
  {SERDES, 4'd13} : path_disable_edge_lane_expected = 1'b0;
  {SAS, 4'd0} : path_disable_edge_lane_expected = 1'b1;
  {SAS, 4'd1} : path_disable_edge_lane_expected = 1'b1;
  {SAS, 4'd2} : path_disable_edge_lane_expected = 1'b1;
  {SAS, 4'd3} : path_disable_edge_lane_expected = 1'b0;
  {SAS, 4'd4} : path_disable_edge_lane_expected = 1'b0;
  {PCIE, 4'd0} : path_disable_edge_lane_expected = 1'b1;
  {PCIE, 4'd1} : path_disable_edge_lane_expected = 1'b1;
  {PCIE, 4'd2} : path_disable_edge_lane_expected = 1'b0;
  {PCIE, 4'd3} : path_disable_edge_lane_expected = 1'b0;
default: path_disable_edge_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : dfe_f1_pol_en_d_lane_expected = 1'b1;
  {USB, 4'd2} : dfe_f1_pol_en_d_lane_expected = 1'b0;
  {SERDES, 4'd0} : dfe_f1_pol_en_d_lane_expected = 1'b1;
  {SERDES, 4'd1} : dfe_f1_pol_en_d_lane_expected = 1'b1;
  {SERDES, 4'd2} : dfe_f1_pol_en_d_lane_expected = 1'b1;
  {SERDES, 4'd3} : dfe_f1_pol_en_d_lane_expected = 1'b1;
  {SERDES, 4'd4} : dfe_f1_pol_en_d_lane_expected = 1'b0;
  {SERDES, 4'd5} : dfe_f1_pol_en_d_lane_expected = 1'b0;
  {SERDES, 4'd6} : dfe_f1_pol_en_d_lane_expected = 1'b0;
  {SERDES, 4'd7} : dfe_f1_pol_en_d_lane_expected = 1'b0;
  {SERDES, 4'd8} : dfe_f1_pol_en_d_lane_expected = 1'b0;
  {SERDES, 4'd9} : dfe_f1_pol_en_d_lane_expected = 1'b0;
  {SERDES, 4'd12} : dfe_f1_pol_en_d_lane_expected = 1'b1;
  {SERDES, 4'd13} : dfe_f1_pol_en_d_lane_expected = 1'b0;
  {SAS, 4'd0} : dfe_f1_pol_en_d_lane_expected = 1'b1;
  {SAS, 4'd1} : dfe_f1_pol_en_d_lane_expected = 1'b1;
  {SAS, 4'd2} : dfe_f1_pol_en_d_lane_expected = 1'b1;
  {SAS, 4'd3} : dfe_f1_pol_en_d_lane_expected = 1'b0;
  {SAS, 4'd4} : dfe_f1_pol_en_d_lane_expected = 1'b0;
  {PCIE, 4'd0} : dfe_f1_pol_en_d_lane_expected = 1'b1;
  {PCIE, 4'd1} : dfe_f1_pol_en_d_lane_expected = 1'b1;
  {PCIE, 4'd2} : dfe_f1_pol_en_d_lane_expected = 1'b0;
  {PCIE, 4'd3} : dfe_f1_pol_en_d_lane_expected = 1'b0;
default: dfe_f1_pol_en_d_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : dfe_f1_pol_en_s_lane_expected = 1'b1;
  {USB, 4'd2} : dfe_f1_pol_en_s_lane_expected = 1'b0;
  {SERDES, 4'd0} : dfe_f1_pol_en_s_lane_expected = 1'b1;
  {SERDES, 4'd1} : dfe_f1_pol_en_s_lane_expected = 1'b1;
  {SERDES, 4'd2} : dfe_f1_pol_en_s_lane_expected = 1'b1;
  {SERDES, 4'd3} : dfe_f1_pol_en_s_lane_expected = 1'b1;
  {SERDES, 4'd4} : dfe_f1_pol_en_s_lane_expected = 1'b0;
  {SERDES, 4'd5} : dfe_f1_pol_en_s_lane_expected = 1'b0;
  {SERDES, 4'd6} : dfe_f1_pol_en_s_lane_expected = 1'b0;
  {SERDES, 4'd7} : dfe_f1_pol_en_s_lane_expected = 1'b0;
  {SERDES, 4'd8} : dfe_f1_pol_en_s_lane_expected = 1'b0;
  {SERDES, 4'd9} : dfe_f1_pol_en_s_lane_expected = 1'b0;
  {SERDES, 4'd12} : dfe_f1_pol_en_s_lane_expected = 1'b1;
  {SERDES, 4'd13} : dfe_f1_pol_en_s_lane_expected = 1'b0;
  {SAS, 4'd0} : dfe_f1_pol_en_s_lane_expected = 1'b1;
  {SAS, 4'd1} : dfe_f1_pol_en_s_lane_expected = 1'b1;
  {SAS, 4'd2} : dfe_f1_pol_en_s_lane_expected = 1'b1;
  {SAS, 4'd3} : dfe_f1_pol_en_s_lane_expected = 1'b0;
  {SAS, 4'd4} : dfe_f1_pol_en_s_lane_expected = 1'b0;
  {PCIE, 4'd0} : dfe_f1_pol_en_s_lane_expected = 1'b1;
  {PCIE, 4'd1} : dfe_f1_pol_en_s_lane_expected = 1'b1;
  {PCIE, 4'd2} : dfe_f1_pol_en_s_lane_expected = 1'b0;
  {PCIE, 4'd3} : dfe_f1_pol_en_s_lane_expected = 1'b0;
default: dfe_f1_pol_en_s_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : dfe_f1_pol_d_lane_expected = 1'b1;
  {USB, 4'd2} : dfe_f1_pol_d_lane_expected = 1'b1;
  {SERDES, 4'd0} : dfe_f1_pol_d_lane_expected = 1'b1;
  {SERDES, 4'd1} : dfe_f1_pol_d_lane_expected = 1'b1;
  {SERDES, 4'd2} : dfe_f1_pol_d_lane_expected = 1'b1;
  {SERDES, 4'd3} : dfe_f1_pol_d_lane_expected = 1'b1;
  {SERDES, 4'd4} : dfe_f1_pol_d_lane_expected = 1'b1;
  {SERDES, 4'd5} : dfe_f1_pol_d_lane_expected = 1'b1;
  {SERDES, 4'd6} : dfe_f1_pol_d_lane_expected = 1'b1;
  {SERDES, 4'd7} : dfe_f1_pol_d_lane_expected = 1'b1;
  {SERDES, 4'd8} : dfe_f1_pol_d_lane_expected = 1'b1;
  {SERDES, 4'd9} : dfe_f1_pol_d_lane_expected = 1'b1;
  {SERDES, 4'd12} : dfe_f1_pol_d_lane_expected = 1'b1;
  {SERDES, 4'd13} : dfe_f1_pol_d_lane_expected = 1'b1;
  {SAS, 4'd0} : dfe_f1_pol_d_lane_expected = 1'b1;
  {SAS, 4'd1} : dfe_f1_pol_d_lane_expected = 1'b1;
  {SAS, 4'd2} : dfe_f1_pol_d_lane_expected = 1'b1;
  {SAS, 4'd3} : dfe_f1_pol_d_lane_expected = 1'b1;
  {SAS, 4'd4} : dfe_f1_pol_d_lane_expected = 1'b1;
  {PCIE, 4'd0} : dfe_f1_pol_d_lane_expected = 1'b1;
  {PCIE, 4'd1} : dfe_f1_pol_d_lane_expected = 1'b1;
  {PCIE, 4'd2} : dfe_f1_pol_d_lane_expected = 1'b1;
  {PCIE, 4'd3} : dfe_f1_pol_d_lane_expected = 1'b1;
default: dfe_f1_pol_d_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : dfe_f1_pol_s_lane_expected = 1'b1;
  {USB, 4'd2} : dfe_f1_pol_s_lane_expected = 1'b1;
  {SERDES, 4'd0} : dfe_f1_pol_s_lane_expected = 1'b1;
  {SERDES, 4'd1} : dfe_f1_pol_s_lane_expected = 1'b1;
  {SERDES, 4'd2} : dfe_f1_pol_s_lane_expected = 1'b1;
  {SERDES, 4'd3} : dfe_f1_pol_s_lane_expected = 1'b1;
  {SERDES, 4'd4} : dfe_f1_pol_s_lane_expected = 1'b1;
  {SERDES, 4'd5} : dfe_f1_pol_s_lane_expected = 1'b1;
  {SERDES, 4'd6} : dfe_f1_pol_s_lane_expected = 1'b1;
  {SERDES, 4'd7} : dfe_f1_pol_s_lane_expected = 1'b1;
  {SERDES, 4'd8} : dfe_f1_pol_s_lane_expected = 1'b1;
  {SERDES, 4'd9} : dfe_f1_pol_s_lane_expected = 1'b1;
  {SERDES, 4'd12} : dfe_f1_pol_s_lane_expected = 1'b1;
  {SERDES, 4'd13} : dfe_f1_pol_s_lane_expected = 1'b1;
  {SAS, 4'd0} : dfe_f1_pol_s_lane_expected = 1'b1;
  {SAS, 4'd1} : dfe_f1_pol_s_lane_expected = 1'b1;
  {SAS, 4'd2} : dfe_f1_pol_s_lane_expected = 1'b1;
  {SAS, 4'd3} : dfe_f1_pol_s_lane_expected = 1'b1;
  {SAS, 4'd4} : dfe_f1_pol_s_lane_expected = 1'b1;
  {PCIE, 4'd0} : dfe_f1_pol_s_lane_expected = 1'b1;
  {PCIE, 4'd1} : dfe_f1_pol_s_lane_expected = 1'b1;
  {PCIE, 4'd2} : dfe_f1_pol_s_lane_expected = 1'b1;
  {PCIE, 4'd3} : dfe_f1_pol_s_lane_expected = 1'b1;
default: dfe_f1_pol_s_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'b1;
  {USB, 4'd2} : reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'b0;
  {SERDES, 4'd0} : reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'b1;
  {SERDES, 4'd1} : reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'b1;
  {SERDES, 4'd2} : reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'b1;
  {SERDES, 4'd3} : reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'b1;
  {SERDES, 4'd4} : reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'b0;
  {SERDES, 4'd5} : reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'b0;
  {SERDES, 4'd6} : reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'b0;
  {SERDES, 4'd7} : reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'b0;
  {SERDES, 4'd8} : reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'b0;
  {SERDES, 4'd9} : reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'b0;
  {SERDES, 4'd12} : reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'b1;
  {SERDES, 4'd13} : reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'b0;
  {SAS, 4'd0} : reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'b1;
  {SAS, 4'd1} : reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'b1;
  {SAS, 4'd2} : reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'b1;
  {SAS, 4'd3} : reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'b0;
  {SAS, 4'd4} : reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'b0;
  {PCIE, 4'd0} : reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'b1;
  {PCIE, 4'd1} : reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'b1;
  {PCIE, 4'd2} : reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'b0;
  {PCIE, 4'd3} : reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'b0;
default: reg_ana_rx_dfe_f1_pol_en_d_force_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'b1;
  {USB, 4'd2} : reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'b0;
  {SERDES, 4'd0} : reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'b1;
  {SERDES, 4'd1} : reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'b1;
  {SERDES, 4'd2} : reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'b1;
  {SERDES, 4'd3} : reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'b1;
  {SERDES, 4'd4} : reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'b0;
  {SERDES, 4'd5} : reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'b0;
  {SERDES, 4'd6} : reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'b0;
  {SERDES, 4'd7} : reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'b0;
  {SERDES, 4'd8} : reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'b0;
  {SERDES, 4'd9} : reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'b0;
  {SERDES, 4'd12} : reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'b1;
  {SERDES, 4'd13} : reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'b0;
  {SAS, 4'd0} : reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'b1;
  {SAS, 4'd1} : reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'b1;
  {SAS, 4'd2} : reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'b1;
  {SAS, 4'd3} : reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'b0;
  {SAS, 4'd4} : reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'b0;
  {PCIE, 4'd0} : reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'b1;
  {PCIE, 4'd1} : reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'b1;
  {PCIE, 4'd2} : reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'b0;
  {PCIE, 4'd3} : reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'b0;
default: reg_ana_rx_dfe_f1_pol_en_s_force_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'b1;
  {USB, 4'd2} : reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'b0;
  {SERDES, 4'd0} : reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'b1;
  {SERDES, 4'd1} : reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'b1;
  {SERDES, 4'd2} : reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'b1;
  {SERDES, 4'd3} : reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'b1;
  {SERDES, 4'd4} : reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'b0;
  {SERDES, 4'd5} : reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'b0;
  {SERDES, 4'd6} : reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'b0;
  {SERDES, 4'd7} : reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'b0;
  {SERDES, 4'd8} : reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'b0;
  {SERDES, 4'd9} : reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'b0;
  {SERDES, 4'd12} : reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'b1;
  {SERDES, 4'd13} : reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'b0;
  {SAS, 4'd0} : reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'b1;
  {SAS, 4'd1} : reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'b1;
  {SAS, 4'd2} : reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'b1;
  {SAS, 4'd3} : reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'b0;
  {SAS, 4'd4} : reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'b0;
  {PCIE, 4'd0} : reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'b1;
  {PCIE, 4'd1} : reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'b1;
  {PCIE, 4'd2} : reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'b0;
  {PCIE, 4'd3} : reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'b0;
default: reg_ana_rx_dfe_f1_pol_d_force_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'b1;
  {USB, 4'd2} : reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'b0;
  {SERDES, 4'd0} : reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'b1;
  {SERDES, 4'd1} : reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'b1;
  {SERDES, 4'd2} : reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'b1;
  {SERDES, 4'd3} : reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'b1;
  {SERDES, 4'd4} : reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'b0;
  {SERDES, 4'd5} : reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'b0;
  {SERDES, 4'd6} : reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'b0;
  {SERDES, 4'd7} : reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'b0;
  {SERDES, 4'd8} : reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'b0;
  {SERDES, 4'd9} : reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'b0;
  {SERDES, 4'd12} : reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'b1;
  {SERDES, 4'd13} : reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'b0;
  {SAS, 4'd0} : reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'b1;
  {SAS, 4'd1} : reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'b1;
  {SAS, 4'd2} : reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'b1;
  {SAS, 4'd3} : reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'b0;
  {SAS, 4'd4} : reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'b0;
  {PCIE, 4'd0} : reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'b1;
  {PCIE, 4'd1} : reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'b1;
  {PCIE, 4'd2} : reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'b0;
  {PCIE, 4'd3} : reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'b0;
default: reg_ana_rx_dfe_f1_pol_s_force_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : reg_dfe_full_rate_mode_lane_expected = 1'b1;
  {USB, 4'd2} : reg_dfe_full_rate_mode_lane_expected = 1'b0;
  {SERDES, 4'd0} : reg_dfe_full_rate_mode_lane_expected = 1'b1;
  {SERDES, 4'd1} : reg_dfe_full_rate_mode_lane_expected = 1'b1;
  {SERDES, 4'd2} : reg_dfe_full_rate_mode_lane_expected = 1'b1;
  {SERDES, 4'd3} : reg_dfe_full_rate_mode_lane_expected = 1'b1;
  {SERDES, 4'd4} : reg_dfe_full_rate_mode_lane_expected = 1'b0;
  {SERDES, 4'd5} : reg_dfe_full_rate_mode_lane_expected = 1'b0;
  {SERDES, 4'd6} : reg_dfe_full_rate_mode_lane_expected = 1'b0;
  {SERDES, 4'd7} : reg_dfe_full_rate_mode_lane_expected = 1'b0;
  {SERDES, 4'd8} : reg_dfe_full_rate_mode_lane_expected = 1'b0;
  {SERDES, 4'd9} : reg_dfe_full_rate_mode_lane_expected = 1'b0;
  {SERDES, 4'd12} : reg_dfe_full_rate_mode_lane_expected = 1'b1;
  {SERDES, 4'd13} : reg_dfe_full_rate_mode_lane_expected = 1'b0;
  {SAS, 4'd0} : reg_dfe_full_rate_mode_lane_expected = 1'b1;
  {SAS, 4'd1} : reg_dfe_full_rate_mode_lane_expected = 1'b1;
  {SAS, 4'd2} : reg_dfe_full_rate_mode_lane_expected = 1'b1;
  {SAS, 4'd3} : reg_dfe_full_rate_mode_lane_expected = 1'b0;
  {SAS, 4'd4} : reg_dfe_full_rate_mode_lane_expected = 1'b0;
  {PCIE, 4'd0} : reg_dfe_full_rate_mode_lane_expected = 1'b1;
  {PCIE, 4'd1} : reg_dfe_full_rate_mode_lane_expected = 1'b1;
  {PCIE, 4'd2} : reg_dfe_full_rate_mode_lane_expected = 1'b0;
  {PCIE, 4'd3} : reg_dfe_full_rate_mode_lane_expected = 1'b0;
default: reg_dfe_full_rate_mode_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : reg_dfe_dis_lane_expected = 1'b0;
  {USB, 4'd2} : reg_dfe_dis_lane_expected = 1'b0;
  {SERDES, 4'd0} : reg_dfe_dis_lane_expected = 1'b1;
  {SERDES, 4'd1} : reg_dfe_dis_lane_expected = 1'b1;
  {SERDES, 4'd2} : reg_dfe_dis_lane_expected = 1'b0;
  {SERDES, 4'd3} : reg_dfe_dis_lane_expected = 1'b0;
  {SERDES, 4'd4} : reg_dfe_dis_lane_expected = 1'b0;
  {SERDES, 4'd5} : reg_dfe_dis_lane_expected = 1'b0;
  {SERDES, 4'd6} : reg_dfe_dis_lane_expected = 1'b0;
  {SERDES, 4'd7} : reg_dfe_dis_lane_expected = 1'b0;
  {SERDES, 4'd8} : reg_dfe_dis_lane_expected = 1'b0;
  {SERDES, 4'd9} : reg_dfe_dis_lane_expected = 1'b0;
  {SERDES, 4'd12} : reg_dfe_dis_lane_expected = 1'b1;
  {SERDES, 4'd13} : reg_dfe_dis_lane_expected = 1'b0;
  {SAS, 4'd0} : reg_dfe_dis_lane_expected = 1'b1;
  {SAS, 4'd1} : reg_dfe_dis_lane_expected = 1'b1;
  {SAS, 4'd2} : reg_dfe_dis_lane_expected = 1'b0;
  {SAS, 4'd3} : reg_dfe_dis_lane_expected = 1'b0;
  {SAS, 4'd4} : reg_dfe_dis_lane_expected = 1'b0;
  {PCIE, 4'd0} : reg_dfe_dis_lane_expected = 1'b1;
  {PCIE, 4'd1} : reg_dfe_dis_lane_expected = 1'b0;
  {PCIE, 4'd2} : reg_dfe_dis_lane_expected = 1'b0;
  {PCIE, 4'd3} : reg_dfe_dis_lane_expected = 1'b0;
default: reg_dfe_dis_lane_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : reg_dfe_tap_settle_scale_lane_expected = 2'b10;
  {USB, 4'd2} : reg_dfe_tap_settle_scale_lane_expected = 2'b01;
  {SERDES, 4'd0} : reg_dfe_tap_settle_scale_lane_expected = 2'b11;
  {SERDES, 4'd1} : reg_dfe_tap_settle_scale_lane_expected = 2'b11;
  {SERDES, 4'd2} : reg_dfe_tap_settle_scale_lane_expected = 2'b10;
  {SERDES, 4'd3} : reg_dfe_tap_settle_scale_lane_expected = 2'b10;
  {SERDES, 4'd4} : reg_dfe_tap_settle_scale_lane_expected = 2'b01;
  {SERDES, 4'd5} : reg_dfe_tap_settle_scale_lane_expected = 2'b01;
  {SERDES, 4'd6} : reg_dfe_tap_settle_scale_lane_expected = 2'b01;
  {SERDES, 4'd7} : reg_dfe_tap_settle_scale_lane_expected = 2'b00;
  {SERDES, 4'd8} : reg_dfe_tap_settle_scale_lane_expected = 2'b00;
  {SERDES, 4'd9} : reg_dfe_tap_settle_scale_lane_expected = 2'b00;
  {SERDES, 4'd12} : reg_dfe_tap_settle_scale_lane_expected = 2'b11;
  {SERDES, 4'd13} : reg_dfe_tap_settle_scale_lane_expected = 2'b00;
  {SAS, 4'd0} : reg_dfe_tap_settle_scale_lane_expected = 2'b11;
  {SAS, 4'd1} : reg_dfe_tap_settle_scale_lane_expected = 2'b11;
  {SAS, 4'd2} : reg_dfe_tap_settle_scale_lane_expected = 2'b10;
  {SAS, 4'd3} : reg_dfe_tap_settle_scale_lane_expected = 2'b01;
  {SAS, 4'd4} : reg_dfe_tap_settle_scale_lane_expected = 2'b00;
  {PCIE, 4'd0} : reg_dfe_tap_settle_scale_lane_expected = 2'b11;
  {PCIE, 4'd1} : reg_dfe_tap_settle_scale_lane_expected = 2'b10;
  {PCIE, 4'd2} : reg_dfe_tap_settle_scale_lane_expected = 2'b01;
  {PCIE, 4'd3} : reg_dfe_tap_settle_scale_lane_expected = 2'b00;
default: reg_dfe_tap_settle_scale_lane_expected = 2'bzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : ffe_data_rate_lane_expected = 4'b0100;
  {USB, 4'd2} : ffe_data_rate_lane_expected = 4'b0110;
  {SERDES, 4'd0} : ffe_data_rate_lane_expected = 4'b0010;
  {SERDES, 4'd1} : ffe_data_rate_lane_expected = 4'b0011;
  {SERDES, 4'd2} : ffe_data_rate_lane_expected = 4'b0100;
  {SERDES, 4'd3} : ffe_data_rate_lane_expected = 4'b0100;
  {SERDES, 4'd4} : ffe_data_rate_lane_expected = 4'b0111;
  {SERDES, 4'd5} : ffe_data_rate_lane_expected = 4'b0111;
  {SERDES, 4'd6} : ffe_data_rate_lane_expected = 4'b0111;
  {SERDES, 4'd7} : ffe_data_rate_lane_expected = 4'b1100;
  {SERDES, 4'd8} : ffe_data_rate_lane_expected = 4'b1101;
  {SERDES, 4'd9} : ffe_data_rate_lane_expected = 4'b1101;
  {SERDES, 4'd12} : ffe_data_rate_lane_expected = 4'b0011;
  {SERDES, 4'd13} : ffe_data_rate_lane_expected = 4'b1011;
  {SAS, 4'd0} : ffe_data_rate_lane_expected = 4'b0010;
  {SAS, 4'd1} : ffe_data_rate_lane_expected = 4'b0011;
  {SAS, 4'd2} : ffe_data_rate_lane_expected = 4'b0100;
  {SAS, 4'd3} : ffe_data_rate_lane_expected = 4'b0111;
  {SAS, 4'd4} : ffe_data_rate_lane_expected = 4'b1011;
  {PCIE, 4'd0} : ffe_data_rate_lane_expected = 4'b0011;
  {PCIE, 4'd1} : ffe_data_rate_lane_expected = 4'b0100;
  {PCIE, 4'd2} : ffe_data_rate_lane_expected = 4'b0101;
  {PCIE, 4'd3} : ffe_data_rate_lane_expected = 4'b1001;
default: ffe_data_rate_lane_expected = 4'bzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : ffe_res1_sel_lane_expected = 4'b0110;
  {USB, 4'd2} : ffe_res1_sel_lane_expected = 4'b0110;
  {SERDES, 4'd0} : ffe_res1_sel_lane_expected = 4'b0110;
  {SERDES, 4'd1} : ffe_res1_sel_lane_expected = 4'b0110;
  {SERDES, 4'd2} : ffe_res1_sel_lane_expected = 4'b0110;
  {SERDES, 4'd3} : ffe_res1_sel_lane_expected = 4'b0110;
  {SERDES, 4'd4} : ffe_res1_sel_lane_expected = 4'b0110;
  {SERDES, 4'd5} : ffe_res1_sel_lane_expected = 4'b0110;
  {SERDES, 4'd6} : ffe_res1_sel_lane_expected = 4'b0110;
  {SERDES, 4'd7} : ffe_res1_sel_lane_expected = 4'b0110;
  {SERDES, 4'd8} : ffe_res1_sel_lane_expected = 4'b0110;
  {SERDES, 4'd9} : ffe_res1_sel_lane_expected = 4'b0110;
  {SERDES, 4'd12} : ffe_res1_sel_lane_expected = 4'b0110;
  {SERDES, 4'd13} : ffe_res1_sel_lane_expected = 4'b0110;
  {SAS, 4'd0} : ffe_res1_sel_lane_expected = 4'b0110;
  {SAS, 4'd1} : ffe_res1_sel_lane_expected = 4'b0110;
  {SAS, 4'd2} : ffe_res1_sel_lane_expected = 4'b0110;
  {SAS, 4'd3} : ffe_res1_sel_lane_expected = 4'b0110;
  {SAS, 4'd4} : ffe_res1_sel_lane_expected = 4'b0110;
  {PCIE, 4'd0} : ffe_res1_sel_lane_expected = 4'b0110;
  {PCIE, 4'd1} : ffe_res1_sel_lane_expected = 4'b0110;
  {PCIE, 4'd2} : ffe_res1_sel_lane_expected = 4'b0110;
  {PCIE, 4'd3} : ffe_res1_sel_lane_expected = 4'b0110;
default: ffe_res1_sel_lane_expected = 4'bzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : ffe_cap1_sel_lane_expected = 4'b1100;
  {USB, 4'd2} : ffe_cap1_sel_lane_expected = 4'b1100;
  {SERDES, 4'd0} : ffe_cap1_sel_lane_expected = 4'b1100;
  {SERDES, 4'd1} : ffe_cap1_sel_lane_expected = 4'b1100;
  {SERDES, 4'd2} : ffe_cap1_sel_lane_expected = 4'b1100;
  {SERDES, 4'd3} : ffe_cap1_sel_lane_expected = 4'b1100;
  {SERDES, 4'd4} : ffe_cap1_sel_lane_expected = 4'b1100;
  {SERDES, 4'd5} : ffe_cap1_sel_lane_expected = 4'b1100;
  {SERDES, 4'd6} : ffe_cap1_sel_lane_expected = 4'b1100;
  {SERDES, 4'd7} : ffe_cap1_sel_lane_expected = 4'b1100;
  {SERDES, 4'd8} : ffe_cap1_sel_lane_expected = 4'b1100;
  {SERDES, 4'd9} : ffe_cap1_sel_lane_expected = 4'b1100;
  {SERDES, 4'd12} : ffe_cap1_sel_lane_expected = 4'b1100;
  {SERDES, 4'd13} : ffe_cap1_sel_lane_expected = 4'b1100;
  {SAS, 4'd0} : ffe_cap1_sel_lane_expected = 4'b1100;
  {SAS, 4'd1} : ffe_cap1_sel_lane_expected = 4'b1100;
  {SAS, 4'd2} : ffe_cap1_sel_lane_expected = 4'b1100;
  {SAS, 4'd3} : ffe_cap1_sel_lane_expected = 4'b1100;
  {SAS, 4'd4} : ffe_cap1_sel_lane_expected = 4'b1100;
  {PCIE, 4'd0} : ffe_cap1_sel_lane_expected = 4'b1100;
  {PCIE, 4'd1} : ffe_cap1_sel_lane_expected = 4'b1100;
  {PCIE, 4'd2} : ffe_cap1_sel_lane_expected = 4'b1100;
  {PCIE, 4'd3} : ffe_cap1_sel_lane_expected = 4'b1100;
default: ffe_cap1_sel_lane_expected = 4'bzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : ffe_res2_sel_e_lane_expected = 4'b0000;
  {USB, 4'd2} : ffe_res2_sel_e_lane_expected = 4'b0000;
  {SERDES, 4'd0} : ffe_res2_sel_e_lane_expected = 4'b0000;
  {SERDES, 4'd1} : ffe_res2_sel_e_lane_expected = 4'b0000;
  {SERDES, 4'd2} : ffe_res2_sel_e_lane_expected = 4'b0000;
  {SERDES, 4'd3} : ffe_res2_sel_e_lane_expected = 4'b0000;
  {SERDES, 4'd4} : ffe_res2_sel_e_lane_expected = 4'b0000;
  {SERDES, 4'd5} : ffe_res2_sel_e_lane_expected = 4'b0000;
  {SERDES, 4'd6} : ffe_res2_sel_e_lane_expected = 4'b0000;
  {SERDES, 4'd7} : ffe_res2_sel_e_lane_expected = 4'b0000;
  {SERDES, 4'd8} : ffe_res2_sel_e_lane_expected = 4'b0000;
  {SERDES, 4'd9} : ffe_res2_sel_e_lane_expected = 4'b0000;
  {SERDES, 4'd12} : ffe_res2_sel_e_lane_expected = 4'b0000;
  {SERDES, 4'd13} : ffe_res2_sel_e_lane_expected = 4'b0000;
  {SAS, 4'd0} : ffe_res2_sel_e_lane_expected = 4'b0000;
  {SAS, 4'd1} : ffe_res2_sel_e_lane_expected = 4'b0000;
  {SAS, 4'd2} : ffe_res2_sel_e_lane_expected = 4'b0000;
  {SAS, 4'd3} : ffe_res2_sel_e_lane_expected = 4'b0000;
  {SAS, 4'd4} : ffe_res2_sel_e_lane_expected = 4'b0000;
  {PCIE, 4'd0} : ffe_res2_sel_e_lane_expected = 4'b0000;
  {PCIE, 4'd1} : ffe_res2_sel_e_lane_expected = 4'b0000;
  {PCIE, 4'd2} : ffe_res2_sel_e_lane_expected = 4'b0000;
  {PCIE, 4'd3} : ffe_res2_sel_e_lane_expected = 4'b0000;
default: ffe_res2_sel_e_lane_expected = 4'bzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : ffe_res2_sel_o_lane_expected = 4'b0000;
  {USB, 4'd2} : ffe_res2_sel_o_lane_expected = 4'b0000;
  {SERDES, 4'd0} : ffe_res2_sel_o_lane_expected = 4'b0000;
  {SERDES, 4'd1} : ffe_res2_sel_o_lane_expected = 4'b0000;
  {SERDES, 4'd2} : ffe_res2_sel_o_lane_expected = 4'b0000;
  {SERDES, 4'd3} : ffe_res2_sel_o_lane_expected = 4'b0000;
  {SERDES, 4'd4} : ffe_res2_sel_o_lane_expected = 4'b0000;
  {SERDES, 4'd5} : ffe_res2_sel_o_lane_expected = 4'b0000;
  {SERDES, 4'd6} : ffe_res2_sel_o_lane_expected = 4'b0000;
  {SERDES, 4'd7} : ffe_res2_sel_o_lane_expected = 4'b0000;
  {SERDES, 4'd8} : ffe_res2_sel_o_lane_expected = 4'b0000;
  {SERDES, 4'd9} : ffe_res2_sel_o_lane_expected = 4'b0000;
  {SERDES, 4'd12} : ffe_res2_sel_o_lane_expected = 4'b0000;
  {SERDES, 4'd13} : ffe_res2_sel_o_lane_expected = 4'b0000;
  {SAS, 4'd0} : ffe_res2_sel_o_lane_expected = 4'b0000;
  {SAS, 4'd1} : ffe_res2_sel_o_lane_expected = 4'b0000;
  {SAS, 4'd2} : ffe_res2_sel_o_lane_expected = 4'b0000;
  {SAS, 4'd3} : ffe_res2_sel_o_lane_expected = 4'b0000;
  {SAS, 4'd4} : ffe_res2_sel_o_lane_expected = 4'b0000;
  {PCIE, 4'd0} : ffe_res2_sel_o_lane_expected = 4'b0000;
  {PCIE, 4'd1} : ffe_res2_sel_o_lane_expected = 4'b0000;
  {PCIE, 4'd2} : ffe_res2_sel_o_lane_expected = 4'b0000;
  {PCIE, 4'd3} : ffe_res2_sel_o_lane_expected = 4'b0000;
default: ffe_res2_sel_o_lane_expected = 4'bzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : ffe_cap2_sel_e_lane_expected = 4'b1111;
  {USB, 4'd2} : ffe_cap2_sel_e_lane_expected = 4'b1111;
  {SERDES, 4'd0} : ffe_cap2_sel_e_lane_expected = 4'b1111;
  {SERDES, 4'd1} : ffe_cap2_sel_e_lane_expected = 4'b1111;
  {SERDES, 4'd2} : ffe_cap2_sel_e_lane_expected = 4'b1111;
  {SERDES, 4'd3} : ffe_cap2_sel_e_lane_expected = 4'b1111;
  {SERDES, 4'd4} : ffe_cap2_sel_e_lane_expected = 4'b1111;
  {SERDES, 4'd5} : ffe_cap2_sel_e_lane_expected = 4'b1111;
  {SERDES, 4'd6} : ffe_cap2_sel_e_lane_expected = 4'b1111;
  {SERDES, 4'd7} : ffe_cap2_sel_e_lane_expected = 4'b1111;
  {SERDES, 4'd8} : ffe_cap2_sel_e_lane_expected = 4'b1111;
  {SERDES, 4'd9} : ffe_cap2_sel_e_lane_expected = 4'b1111;
  {SERDES, 4'd12} : ffe_cap2_sel_e_lane_expected = 4'b1111;
  {SERDES, 4'd13} : ffe_cap2_sel_e_lane_expected = 4'b1111;
  {SAS, 4'd0} : ffe_cap2_sel_e_lane_expected = 4'b1111;
  {SAS, 4'd1} : ffe_cap2_sel_e_lane_expected = 4'b1111;
  {SAS, 4'd2} : ffe_cap2_sel_e_lane_expected = 4'b1111;
  {SAS, 4'd3} : ffe_cap2_sel_e_lane_expected = 4'b1111;
  {SAS, 4'd4} : ffe_cap2_sel_e_lane_expected = 4'b1111;
  {PCIE, 4'd0} : ffe_cap2_sel_e_lane_expected = 4'b1111;
  {PCIE, 4'd1} : ffe_cap2_sel_e_lane_expected = 4'b1111;
  {PCIE, 4'd2} : ffe_cap2_sel_e_lane_expected = 4'b1111;
  {PCIE, 4'd3} : ffe_cap2_sel_e_lane_expected = 4'b1111;
default: ffe_cap2_sel_e_lane_expected = 4'bzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : ffe_cap2_sel_o_lane_expected = 4'b1111;
  {USB, 4'd2} : ffe_cap2_sel_o_lane_expected = 4'b1111;
  {SERDES, 4'd0} : ffe_cap2_sel_o_lane_expected = 4'b1111;
  {SERDES, 4'd1} : ffe_cap2_sel_o_lane_expected = 4'b1111;
  {SERDES, 4'd2} : ffe_cap2_sel_o_lane_expected = 4'b1111;
  {SERDES, 4'd3} : ffe_cap2_sel_o_lane_expected = 4'b1111;
  {SERDES, 4'd4} : ffe_cap2_sel_o_lane_expected = 4'b1111;
  {SERDES, 4'd5} : ffe_cap2_sel_o_lane_expected = 4'b1111;
  {SERDES, 4'd6} : ffe_cap2_sel_o_lane_expected = 4'b1111;
  {SERDES, 4'd7} : ffe_cap2_sel_o_lane_expected = 4'b1111;
  {SERDES, 4'd8} : ffe_cap2_sel_o_lane_expected = 4'b1111;
  {SERDES, 4'd9} : ffe_cap2_sel_o_lane_expected = 4'b1111;
  {SERDES, 4'd12} : ffe_cap2_sel_o_lane_expected = 4'b1111;
  {SERDES, 4'd13} : ffe_cap2_sel_o_lane_expected = 4'b1111;
  {SAS, 4'd0} : ffe_cap2_sel_o_lane_expected = 4'b1111;
  {SAS, 4'd1} : ffe_cap2_sel_o_lane_expected = 4'b1111;
  {SAS, 4'd2} : ffe_cap2_sel_o_lane_expected = 4'b1111;
  {SAS, 4'd3} : ffe_cap2_sel_o_lane_expected = 4'b1111;
  {SAS, 4'd4} : ffe_cap2_sel_o_lane_expected = 4'b1111;
  {PCIE, 4'd0} : ffe_cap2_sel_o_lane_expected = 4'b1111;
  {PCIE, 4'd1} : ffe_cap2_sel_o_lane_expected = 4'b1111;
  {PCIE, 4'd2} : ffe_cap2_sel_o_lane_expected = 4'b1111;
  {PCIE, 4'd3} : ffe_cap2_sel_o_lane_expected = 4'b1111;
default: ffe_cap2_sel_o_lane_expected = 4'bzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : rxdll_temp_a_lane_expected = 8'b00011011;
  {USB, 4'd2} : rxdll_temp_a_lane_expected = 8'b00011011;
  {SERDES, 4'd0} : rxdll_temp_a_lane_expected = 8'b00011011;
  {SERDES, 4'd1} : rxdll_temp_a_lane_expected = 8'b00100001;
  {SERDES, 4'd2} : rxdll_temp_a_lane_expected = 8'b00011011;
  {SERDES, 4'd3} : rxdll_temp_a_lane_expected = 8'b00100001;
  {SERDES, 4'd4} : rxdll_temp_a_lane_expected = 8'b00011011;
  {SERDES, 4'd5} : rxdll_temp_a_lane_expected = 8'b00100001;
  {SERDES, 4'd6} : rxdll_temp_a_lane_expected = 8'b00100001;
  {SERDES, 4'd7} : rxdll_temp_a_lane_expected = 8'b00100001;
  {SERDES, 4'd8} : rxdll_temp_a_lane_expected = 8'b00100100;
  {SERDES, 4'd9} : rxdll_temp_a_lane_expected = 8'b00100100;
  {SERDES, 4'd12} : rxdll_temp_a_lane_expected = 8'b00011011;
  {SERDES, 4'd13} : rxdll_temp_a_lane_expected = 8'b00011011;
  {SAS, 4'd0} : rxdll_temp_a_lane_expected = 8'b00100001;
  {SAS, 4'd1} : rxdll_temp_a_lane_expected = 8'b00100001;
  {SAS, 4'd2} : rxdll_temp_a_lane_expected = 8'b00100001;
  {SAS, 4'd3} : rxdll_temp_a_lane_expected = 8'b00100001;
  {SAS, 4'd4} : rxdll_temp_a_lane_expected = 8'b00011011;
  {PCIE, 4'd0} : rxdll_temp_a_lane_expected = 8'b00011011;
  {PCIE, 4'd1} : rxdll_temp_a_lane_expected = 8'b00011011;
  {PCIE, 4'd2} : rxdll_temp_a_lane_expected = 8'b00011110;
  {PCIE, 4'd3} : rxdll_temp_a_lane_expected = 8'b00011110;
default: rxdll_temp_a_lane_expected = 8'bzzzzzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0])
case ( {phy_mode_bit[2:0], gen[3:0]} )
  {USB, 4'd1} : rxdll_temp_b_lane_expected = 8'b10100000;
  {USB, 4'd2} : rxdll_temp_b_lane_expected = 8'b10100000;
  {SERDES, 4'd0} : rxdll_temp_b_lane_expected = 8'b10100000;
  {SERDES, 4'd1} : rxdll_temp_b_lane_expected = 8'b10100000;
  {SERDES, 4'd2} : rxdll_temp_b_lane_expected = 8'b10100000;
  {SERDES, 4'd3} : rxdll_temp_b_lane_expected = 8'b10100000;
  {SERDES, 4'd4} : rxdll_temp_b_lane_expected = 8'b10100000;
  {SERDES, 4'd5} : rxdll_temp_b_lane_expected = 8'b10100000;
  {SERDES, 4'd6} : rxdll_temp_b_lane_expected = 8'b10100000;
  {SERDES, 4'd7} : rxdll_temp_b_lane_expected = 8'b10100000;
  {SERDES, 4'd8} : rxdll_temp_b_lane_expected = 8'b10101100;
  {SERDES, 4'd9} : rxdll_temp_b_lane_expected = 8'b10101100;
  {SERDES, 4'd12} : rxdll_temp_b_lane_expected = 8'b10100000;
  {SERDES, 4'd13} : rxdll_temp_b_lane_expected = 8'b10100000;
  {SAS, 4'd0} : rxdll_temp_b_lane_expected = 8'b10100000;
  {SAS, 4'd1} : rxdll_temp_b_lane_expected = 8'b10100000;
  {SAS, 4'd2} : rxdll_temp_b_lane_expected = 8'b10100000;
  {SAS, 4'd3} : rxdll_temp_b_lane_expected = 8'b10100000;
  {SAS, 4'd4} : rxdll_temp_b_lane_expected = 8'b10100000;
  {PCIE, 4'd0} : rxdll_temp_b_lane_expected = 8'b10100000;
  {PCIE, 4'd1} : rxdll_temp_b_lane_expected = 8'b10100000;
  {PCIE, 4'd2} : rxdll_temp_b_lane_expected = 8'b10100000;
  {PCIE, 4'd3} : rxdll_temp_b_lane_expected = 8'b10100000;
default: rxdll_temp_b_lane_expected = 8'bzzzzzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel} )
  {USB, 4'd1, 5'd0, 1'd0} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd1, 5'd1, 1'd0} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd1, 5'd2, 1'd0} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd1, 5'd3, 1'd0} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd1, 5'd4, 1'd0} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd1, 5'd5, 1'd0} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd1, 5'd6, 1'd0} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd1, 5'd7, 1'd0} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd2, 5'd0, 1'd0} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd2, 5'd1, 1'd0} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd2, 5'd2, 1'd0} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd2, 5'd3, 1'd0} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd2, 5'd4, 1'd0} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd2, 5'd5, 1'd0} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd2, 5'd6, 1'd0} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd2, 5'd7, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd0, 5'd0, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd0, 5'd1, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd0, 5'd2, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd0, 5'd3, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd0, 5'd4, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd0, 5'd5, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd0, 5'd6, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd0, 5'd7, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd1, 5'd0, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd1, 5'd1, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd1, 5'd2, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd1, 5'd3, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd1, 5'd4, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd1, 5'd5, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd1, 5'd6, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd1, 5'd7, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd2, 5'd0, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd2, 5'd1, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd2, 5'd2, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd2, 5'd3, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd2, 5'd4, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd2, 5'd5, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd2, 5'd6, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd2, 5'd7, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd3, 5'd0, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd3, 5'd1, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd3, 5'd2, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd3, 5'd3, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd3, 5'd4, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd3, 5'd5, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd3, 5'd6, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd3, 5'd7, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd4, 5'd0, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd4, 5'd1, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd4, 5'd2, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd4, 5'd3, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd4, 5'd4, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd4, 5'd5, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd4, 5'd6, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd4, 5'd7, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd5, 5'd0, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd5, 5'd1, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd5, 5'd2, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd5, 5'd3, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd5, 5'd4, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd5, 5'd5, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd5, 5'd6, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd5, 5'd7, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd6, 5'd0, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd6, 5'd1, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd6, 5'd2, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd6, 5'd3, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd6, 5'd4, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd6, 5'd5, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd6, 5'd6, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd6, 5'd7, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd7, 5'd0, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd7, 5'd1, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd7, 5'd2, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd7, 5'd3, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd7, 5'd4, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd7, 5'd5, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd7, 5'd6, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd7, 5'd7, 1'd0} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd8, 5'd0, 1'd0} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd8, 5'd1, 1'd0} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd8, 5'd2, 1'd0} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd8, 5'd3, 1'd0} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd8, 5'd4, 1'd0} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd8, 5'd5, 1'd0} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd8, 5'd6, 1'd0} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd8, 5'd7, 1'd0} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd9, 5'd0, 1'd0} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd9, 5'd1, 1'd0} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd9, 5'd2, 1'd0} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd9, 5'd3, 1'd0} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd9, 5'd4, 1'd0} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd9, 5'd5, 1'd0} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd9, 5'd6, 1'd0} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd9, 5'd7, 1'd0} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd12, 5'd0, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd12, 5'd1, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd12, 5'd2, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd12, 5'd3, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd12, 5'd4, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd12, 5'd5, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd12, 5'd6, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd12, 5'd7, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd13, 5'd0, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd13, 5'd1, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd13, 5'd2, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd13, 5'd3, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd13, 5'd4, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd13, 5'd5, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd13, 5'd6, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd13, 5'd7, 1'd0} : pll_reg_sel_expected = 3'b000;
  {SAS, 4'd0, 5'd0, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd0, 5'd1, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd0, 5'd2, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd0, 5'd3, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd0, 5'd4, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd0, 5'd5, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd0, 5'd6, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd0, 5'd7, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd1, 5'd0, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd1, 5'd1, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd1, 5'd2, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd1, 5'd3, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd1, 5'd4, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd1, 5'd5, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd1, 5'd6, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd1, 5'd7, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd2, 5'd0, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd2, 5'd1, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd2, 5'd2, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd2, 5'd3, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd2, 5'd4, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd2, 5'd5, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd2, 5'd6, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd2, 5'd7, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd3, 5'd0, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd3, 5'd1, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd3, 5'd2, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd3, 5'd3, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd3, 5'd4, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd3, 5'd5, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd3, 5'd6, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd3, 5'd7, 1'd0} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd4, 5'd0, 1'd0} : pll_reg_sel_expected = 3'b001;
  {SAS, 4'd4, 5'd1, 1'd0} : pll_reg_sel_expected = 3'b001;
  {SAS, 4'd4, 5'd2, 1'd0} : pll_reg_sel_expected = 3'b001;
  {SAS, 4'd4, 5'd3, 1'd0} : pll_reg_sel_expected = 3'b001;
  {SAS, 4'd4, 5'd4, 1'd0} : pll_reg_sel_expected = 3'b001;
  {SAS, 4'd4, 5'd5, 1'd0} : pll_reg_sel_expected = 3'b001;
  {SAS, 4'd4, 5'd6, 1'd0} : pll_reg_sel_expected = 3'b001;
  {SAS, 4'd4, 5'd7, 1'd0} : pll_reg_sel_expected = 3'b001;
  {PCIE, 4'd2, 5'd0, 1'd0} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd2, 5'd1, 1'd0} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd2, 5'd2, 1'd0} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd2, 5'd3, 1'd0} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd2, 5'd4, 1'd0} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd2, 5'd5, 1'd0} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd2, 5'd6, 1'd0} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd2, 5'd7, 1'd0} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd3, 5'd0, 1'd0} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd3, 5'd1, 1'd0} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd3, 5'd2, 1'd0} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd3, 5'd3, 1'd0} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd3, 5'd4, 1'd0} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd3, 5'd5, 1'd0} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd3, 5'd6, 1'd0} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd3, 5'd7, 1'd0} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd1, 5'd0, 1'd1} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd1, 5'd1, 1'd1} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd1, 5'd2, 1'd1} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd1, 5'd3, 1'd1} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd1, 5'd4, 1'd1} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd1, 5'd5, 1'd1} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd1, 5'd6, 1'd1} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd1, 5'd7, 1'd1} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd2, 5'd0, 1'd1} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd2, 5'd1, 1'd1} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd2, 5'd2, 1'd1} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd2, 5'd3, 1'd1} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd2, 5'd4, 1'd1} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd2, 5'd5, 1'd1} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd2, 5'd6, 1'd1} : pll_reg_sel_expected = 3'b000;
  {USB, 4'd2, 5'd7, 1'd1} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd0, 5'd0, 1'd1} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd0, 5'd1, 1'd1} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd0, 5'd2, 1'd1} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd0, 5'd3, 1'd1} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd0, 5'd4, 1'd1} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd0, 5'd5, 1'd1} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd0, 5'd6, 1'd1} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd0, 5'd7, 1'd1} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd1, 5'd0, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd1, 5'd1, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd1, 5'd2, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd1, 5'd3, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd1, 5'd4, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd1, 5'd5, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd1, 5'd6, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd1, 5'd7, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd2, 5'd0, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd2, 5'd1, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd2, 5'd2, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd2, 5'd3, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd2, 5'd4, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd2, 5'd5, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd2, 5'd6, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd2, 5'd7, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd3, 5'd0, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd3, 5'd1, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd3, 5'd2, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd3, 5'd3, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd3, 5'd4, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd3, 5'd5, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd3, 5'd6, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd3, 5'd7, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd4, 5'd0, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd4, 5'd1, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd4, 5'd2, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd4, 5'd3, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd4, 5'd4, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd4, 5'd5, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd4, 5'd6, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd4, 5'd7, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd5, 5'd0, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd5, 5'd1, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd5, 5'd2, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd5, 5'd3, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd5, 5'd4, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd5, 5'd5, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd5, 5'd6, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd5, 5'd7, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd6, 5'd0, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd6, 5'd1, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd6, 5'd2, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd6, 5'd3, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd6, 5'd4, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd6, 5'd5, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd6, 5'd6, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd6, 5'd7, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd7, 5'd0, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd7, 5'd1, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd7, 5'd2, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd7, 5'd3, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd7, 5'd4, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd7, 5'd5, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd7, 5'd6, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd7, 5'd7, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd8, 5'd0, 1'd1} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd8, 5'd1, 1'd1} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd8, 5'd2, 1'd1} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd8, 5'd3, 1'd1} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd8, 5'd4, 1'd1} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd8, 5'd5, 1'd1} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd8, 5'd6, 1'd1} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd8, 5'd7, 1'd1} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd9, 5'd0, 1'd1} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd9, 5'd1, 1'd1} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd9, 5'd2, 1'd1} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd9, 5'd3, 1'd1} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd9, 5'd4, 1'd1} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd9, 5'd5, 1'd1} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd9, 5'd6, 1'd1} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd9, 5'd7, 1'd1} : pll_reg_sel_expected = 3'b100;
  {SERDES, 4'd12, 5'd0, 1'd1} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd12, 5'd1, 1'd1} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd12, 5'd2, 1'd1} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd12, 5'd3, 1'd1} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd12, 5'd4, 1'd1} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd12, 5'd5, 1'd1} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd12, 5'd6, 1'd1} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd12, 5'd7, 1'd1} : pll_reg_sel_expected = 3'b000;
  {SERDES, 4'd13, 5'd0, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd13, 5'd1, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd13, 5'd2, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd13, 5'd3, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd13, 5'd4, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd13, 5'd5, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd13, 5'd6, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SERDES, 4'd13, 5'd7, 1'd1} : pll_reg_sel_expected = 3'b011;
  {SAS, 4'd0, 5'd0, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd0, 5'd1, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd0, 5'd2, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd0, 5'd3, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd0, 5'd4, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd0, 5'd5, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd0, 5'd6, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd0, 5'd7, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd1, 5'd0, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd1, 5'd1, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd1, 5'd2, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd1, 5'd3, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd1, 5'd4, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd1, 5'd5, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd1, 5'd6, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd1, 5'd7, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd2, 5'd0, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd2, 5'd1, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd2, 5'd2, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd2, 5'd3, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd2, 5'd4, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd2, 5'd5, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd2, 5'd6, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd2, 5'd7, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd3, 5'd0, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd3, 5'd1, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd3, 5'd2, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd3, 5'd3, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd3, 5'd4, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd3, 5'd5, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd3, 5'd6, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd3, 5'd7, 1'd1} : pll_reg_sel_expected = 3'b010;
  {SAS, 4'd4, 5'd0, 1'd1} : pll_reg_sel_expected = 3'b001;
  {SAS, 4'd4, 5'd1, 1'd1} : pll_reg_sel_expected = 3'b001;
  {SAS, 4'd4, 5'd2, 1'd1} : pll_reg_sel_expected = 3'b001;
  {SAS, 4'd4, 5'd3, 1'd1} : pll_reg_sel_expected = 3'b001;
  {SAS, 4'd4, 5'd4, 1'd1} : pll_reg_sel_expected = 3'b001;
  {SAS, 4'd4, 5'd5, 1'd1} : pll_reg_sel_expected = 3'b001;
  {SAS, 4'd4, 5'd6, 1'd1} : pll_reg_sel_expected = 3'b001;
  {SAS, 4'd4, 5'd7, 1'd1} : pll_reg_sel_expected = 3'b001;
  {PCIE, 4'd2, 5'd0, 1'd1} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd2, 5'd1, 1'd1} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd2, 5'd2, 1'd1} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd2, 5'd3, 1'd1} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd2, 5'd4, 1'd1} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd2, 5'd5, 1'd1} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd2, 5'd6, 1'd1} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd2, 5'd7, 1'd1} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd3, 5'd0, 1'd1} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd3, 5'd1, 1'd1} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd3, 5'd2, 1'd1} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd3, 5'd3, 1'd1} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd3, 5'd4, 1'd1} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd3, 5'd5, 1'd1} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd3, 5'd6, 1'd1} : pll_reg_sel_expected = 3'b000;
  {PCIE, 4'd3, 5'd7, 1'd1} : pll_reg_sel_expected = 3'b000;
default: pll_reg_sel_expected = 3'bzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel} )
  {USB, 4'd1, 5'd0, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd1, 5'd1, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd1, 5'd2, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd1, 5'd3, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd1, 5'd4, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd1, 5'd5, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd1, 5'd6, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd1, 5'd7, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd2, 5'd0, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd2, 5'd1, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd2, 5'd2, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd2, 5'd3, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd2, 5'd4, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd2, 5'd5, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd2, 5'd6, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd2, 5'd7, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd0, 5'd0, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd0, 5'd1, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd0, 5'd2, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd0, 5'd3, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd0, 5'd4, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd0, 5'd5, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd0, 5'd6, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd0, 5'd7, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd1, 5'd0, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd1, 5'd1, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd1, 5'd2, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd1, 5'd3, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd1, 5'd4, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd1, 5'd5, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd1, 5'd6, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd1, 5'd7, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd2, 5'd0, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd2, 5'd1, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd2, 5'd2, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd2, 5'd3, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd2, 5'd4, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd2, 5'd5, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd2, 5'd6, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd2, 5'd7, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd3, 5'd0, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd3, 5'd1, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd3, 5'd2, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd3, 5'd3, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd3, 5'd4, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd3, 5'd5, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd3, 5'd6, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd3, 5'd7, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd4, 5'd0, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd4, 5'd1, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd4, 5'd2, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd4, 5'd3, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd4, 5'd4, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd4, 5'd5, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd4, 5'd6, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd4, 5'd7, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd5, 5'd0, 1'd0} : pll_rate_sel_expected = 4'b0010;
  {SERDES, 4'd5, 5'd1, 1'd0} : pll_rate_sel_expected = 4'b0010;
  {SERDES, 4'd5, 5'd2, 1'd0} : pll_rate_sel_expected = 4'b0010;
  {SERDES, 4'd5, 5'd3, 1'd0} : pll_rate_sel_expected = 4'b0010;
  {SERDES, 4'd5, 5'd4, 1'd0} : pll_rate_sel_expected = 4'b0010;
  {SERDES, 4'd5, 5'd5, 1'd0} : pll_rate_sel_expected = 4'b0010;
  {SERDES, 4'd5, 5'd6, 1'd0} : pll_rate_sel_expected = 4'b0010;
  {SERDES, 4'd5, 5'd7, 1'd0} : pll_rate_sel_expected = 4'b0010;
  {SERDES, 4'd6, 5'd0, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd6, 5'd1, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd6, 5'd2, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd6, 5'd3, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd6, 5'd4, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd6, 5'd5, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd6, 5'd6, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd6, 5'd7, 1'd0} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd7, 5'd0, 1'd0} : pll_rate_sel_expected = 4'b0100;
  {SERDES, 4'd7, 5'd1, 1'd0} : pll_rate_sel_expected = 4'b0100;
  {SERDES, 4'd7, 5'd2, 1'd0} : pll_rate_sel_expected = 4'b0100;
  {SERDES, 4'd7, 5'd3, 1'd0} : pll_rate_sel_expected = 4'b0100;
  {SERDES, 4'd7, 5'd4, 1'd0} : pll_rate_sel_expected = 4'b0100;
  {SERDES, 4'd7, 5'd5, 1'd0} : pll_rate_sel_expected = 4'b0100;
  {SERDES, 4'd7, 5'd6, 1'd0} : pll_rate_sel_expected = 4'b0100;
  {SERDES, 4'd7, 5'd7, 1'd0} : pll_rate_sel_expected = 4'b0100;
  {SERDES, 4'd8, 5'd0, 1'd0} : pll_rate_sel_expected = 4'b0101;
  {SERDES, 4'd8, 5'd1, 1'd0} : pll_rate_sel_expected = 4'b0101;
  {SERDES, 4'd8, 5'd2, 1'd0} : pll_rate_sel_expected = 4'b0101;
  {SERDES, 4'd8, 5'd3, 1'd0} : pll_rate_sel_expected = 4'b0101;
  {SERDES, 4'd8, 5'd4, 1'd0} : pll_rate_sel_expected = 4'b0101;
  {SERDES, 4'd8, 5'd5, 1'd0} : pll_rate_sel_expected = 4'b0101;
  {SERDES, 4'd8, 5'd6, 1'd0} : pll_rate_sel_expected = 4'b0101;
  {SERDES, 4'd8, 5'd7, 1'd0} : pll_rate_sel_expected = 4'b0101;
  {SERDES, 4'd9, 5'd0, 1'd0} : pll_rate_sel_expected = 4'b0110;
  {SERDES, 4'd9, 5'd1, 1'd0} : pll_rate_sel_expected = 4'b0110;
  {SERDES, 4'd9, 5'd2, 1'd0} : pll_rate_sel_expected = 4'b0110;
  {SERDES, 4'd9, 5'd3, 1'd0} : pll_rate_sel_expected = 4'b0110;
  {SERDES, 4'd9, 5'd4, 1'd0} : pll_rate_sel_expected = 4'b0110;
  {SERDES, 4'd9, 5'd5, 1'd0} : pll_rate_sel_expected = 4'b0110;
  {SERDES, 4'd9, 5'd6, 1'd0} : pll_rate_sel_expected = 4'b0110;
  {SERDES, 4'd9, 5'd7, 1'd0} : pll_rate_sel_expected = 4'b0110;
  {SERDES, 4'd12, 5'd0, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd12, 5'd1, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd12, 5'd2, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd12, 5'd3, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd12, 5'd4, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd12, 5'd5, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd12, 5'd6, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd12, 5'd7, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd13, 5'd0, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd13, 5'd1, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd13, 5'd2, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd13, 5'd3, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd13, 5'd4, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd13, 5'd5, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd13, 5'd6, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd13, 5'd7, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd0, 5'd0, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd0, 5'd1, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd0, 5'd2, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd0, 5'd3, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd0, 5'd4, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd0, 5'd5, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd0, 5'd6, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd0, 5'd7, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd1, 5'd0, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd1, 5'd1, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd1, 5'd2, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd1, 5'd3, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd1, 5'd4, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd1, 5'd5, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd1, 5'd6, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd1, 5'd7, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd2, 5'd0, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd2, 5'd1, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd2, 5'd2, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd2, 5'd3, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd2, 5'd4, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd2, 5'd5, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd2, 5'd6, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd2, 5'd7, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd3, 5'd0, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd3, 5'd1, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd3, 5'd2, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd3, 5'd3, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd3, 5'd4, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd3, 5'd5, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd3, 5'd6, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd3, 5'd7, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd4, 5'd0, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SAS, 4'd4, 5'd1, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SAS, 4'd4, 5'd2, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SAS, 4'd4, 5'd3, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SAS, 4'd4, 5'd4, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SAS, 4'd4, 5'd5, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SAS, 4'd4, 5'd6, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {SAS, 4'd4, 5'd7, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd0, 5'd0, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd0, 5'd1, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd0, 5'd2, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd0, 5'd3, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd0, 5'd4, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd0, 5'd5, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd0, 5'd6, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd0, 5'd7, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd1, 5'd0, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd1, 5'd1, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd1, 5'd2, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd1, 5'd3, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd1, 5'd4, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd1, 5'd5, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd1, 5'd6, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd1, 5'd7, 1'd0} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd2, 5'd0, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd2, 5'd1, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd2, 5'd2, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd2, 5'd3, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd2, 5'd4, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd2, 5'd5, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd2, 5'd6, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd2, 5'd7, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd3, 5'd0, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd3, 5'd1, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd3, 5'd2, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd3, 5'd3, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd3, 5'd4, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd3, 5'd5, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd3, 5'd6, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd3, 5'd7, 1'd0} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd1, 5'd0, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd1, 5'd1, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd1, 5'd2, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd1, 5'd3, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd1, 5'd4, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd1, 5'd5, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd1, 5'd6, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd1, 5'd7, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd2, 5'd0, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd2, 5'd1, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd2, 5'd2, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd2, 5'd3, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd2, 5'd4, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd2, 5'd5, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd2, 5'd6, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {USB, 4'd2, 5'd7, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd0, 5'd0, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd0, 5'd1, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd0, 5'd2, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd0, 5'd3, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd0, 5'd4, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd0, 5'd5, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd0, 5'd6, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd0, 5'd7, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd1, 5'd0, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd1, 5'd1, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd1, 5'd2, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd1, 5'd3, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd1, 5'd4, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd1, 5'd5, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd1, 5'd6, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd1, 5'd7, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd2, 5'd0, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd2, 5'd1, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd2, 5'd2, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd2, 5'd3, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd2, 5'd4, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd2, 5'd5, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd2, 5'd6, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd2, 5'd7, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd3, 5'd0, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd3, 5'd1, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd3, 5'd2, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd3, 5'd3, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd3, 5'd4, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd3, 5'd5, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd3, 5'd6, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd3, 5'd7, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd4, 5'd0, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd4, 5'd1, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd4, 5'd2, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd4, 5'd3, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd4, 5'd4, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd4, 5'd5, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd4, 5'd6, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd4, 5'd7, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd5, 5'd0, 1'd1} : pll_rate_sel_expected = 4'b0010;
  {SERDES, 4'd5, 5'd1, 1'd1} : pll_rate_sel_expected = 4'b0010;
  {SERDES, 4'd5, 5'd2, 1'd1} : pll_rate_sel_expected = 4'b0010;
  {SERDES, 4'd5, 5'd3, 1'd1} : pll_rate_sel_expected = 4'b0010;
  {SERDES, 4'd5, 5'd4, 1'd1} : pll_rate_sel_expected = 4'b0010;
  {SERDES, 4'd5, 5'd5, 1'd1} : pll_rate_sel_expected = 4'b0010;
  {SERDES, 4'd5, 5'd6, 1'd1} : pll_rate_sel_expected = 4'b0010;
  {SERDES, 4'd5, 5'd7, 1'd1} : pll_rate_sel_expected = 4'b0010;
  {SERDES, 4'd6, 5'd0, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd6, 5'd1, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd6, 5'd2, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd6, 5'd3, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd6, 5'd4, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd6, 5'd5, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd6, 5'd6, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd6, 5'd7, 1'd1} : pll_rate_sel_expected = 4'b0011;
  {SERDES, 4'd7, 5'd0, 1'd1} : pll_rate_sel_expected = 4'b0100;
  {SERDES, 4'd7, 5'd1, 1'd1} : pll_rate_sel_expected = 4'b0100;
  {SERDES, 4'd7, 5'd2, 1'd1} : pll_rate_sel_expected = 4'b0100;
  {SERDES, 4'd7, 5'd3, 1'd1} : pll_rate_sel_expected = 4'b0100;
  {SERDES, 4'd7, 5'd4, 1'd1} : pll_rate_sel_expected = 4'b0100;
  {SERDES, 4'd7, 5'd5, 1'd1} : pll_rate_sel_expected = 4'b0100;
  {SERDES, 4'd7, 5'd6, 1'd1} : pll_rate_sel_expected = 4'b0100;
  {SERDES, 4'd7, 5'd7, 1'd1} : pll_rate_sel_expected = 4'b0100;
  {SERDES, 4'd8, 5'd0, 1'd1} : pll_rate_sel_expected = 4'b0101;
  {SERDES, 4'd8, 5'd1, 1'd1} : pll_rate_sel_expected = 4'b0101;
  {SERDES, 4'd8, 5'd2, 1'd1} : pll_rate_sel_expected = 4'b0101;
  {SERDES, 4'd8, 5'd3, 1'd1} : pll_rate_sel_expected = 4'b0101;
  {SERDES, 4'd8, 5'd4, 1'd1} : pll_rate_sel_expected = 4'b0101;
  {SERDES, 4'd8, 5'd5, 1'd1} : pll_rate_sel_expected = 4'b0101;
  {SERDES, 4'd8, 5'd6, 1'd1} : pll_rate_sel_expected = 4'b0101;
  {SERDES, 4'd8, 5'd7, 1'd1} : pll_rate_sel_expected = 4'b0101;
  {SERDES, 4'd9, 5'd0, 1'd1} : pll_rate_sel_expected = 4'b0110;
  {SERDES, 4'd9, 5'd1, 1'd1} : pll_rate_sel_expected = 4'b0110;
  {SERDES, 4'd9, 5'd2, 1'd1} : pll_rate_sel_expected = 4'b0110;
  {SERDES, 4'd9, 5'd3, 1'd1} : pll_rate_sel_expected = 4'b0110;
  {SERDES, 4'd9, 5'd4, 1'd1} : pll_rate_sel_expected = 4'b0110;
  {SERDES, 4'd9, 5'd5, 1'd1} : pll_rate_sel_expected = 4'b0110;
  {SERDES, 4'd9, 5'd6, 1'd1} : pll_rate_sel_expected = 4'b0110;
  {SERDES, 4'd9, 5'd7, 1'd1} : pll_rate_sel_expected = 4'b0110;
  {SERDES, 4'd12, 5'd0, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd12, 5'd1, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd12, 5'd2, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd12, 5'd3, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd12, 5'd4, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd12, 5'd5, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd12, 5'd6, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd12, 5'd7, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SERDES, 4'd13, 5'd0, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd13, 5'd1, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd13, 5'd2, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd13, 5'd3, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd13, 5'd4, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd13, 5'd5, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd13, 5'd6, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SERDES, 4'd13, 5'd7, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd0, 5'd0, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd0, 5'd1, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd0, 5'd2, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd0, 5'd3, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd0, 5'd4, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd0, 5'd5, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd0, 5'd6, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd0, 5'd7, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd1, 5'd0, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd1, 5'd1, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd1, 5'd2, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd1, 5'd3, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd1, 5'd4, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd1, 5'd5, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd1, 5'd6, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd1, 5'd7, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd2, 5'd0, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd2, 5'd1, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd2, 5'd2, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd2, 5'd3, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd2, 5'd4, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd2, 5'd5, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd2, 5'd6, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd2, 5'd7, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd3, 5'd0, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd3, 5'd1, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd3, 5'd2, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd3, 5'd3, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd3, 5'd4, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd3, 5'd5, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd3, 5'd6, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd3, 5'd7, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {SAS, 4'd4, 5'd0, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SAS, 4'd4, 5'd1, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SAS, 4'd4, 5'd2, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SAS, 4'd4, 5'd3, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SAS, 4'd4, 5'd4, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SAS, 4'd4, 5'd5, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SAS, 4'd4, 5'd6, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {SAS, 4'd4, 5'd7, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd0, 5'd0, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd0, 5'd1, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd0, 5'd2, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd0, 5'd3, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd0, 5'd4, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd0, 5'd5, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd0, 5'd6, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd0, 5'd7, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd1, 5'd0, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd1, 5'd1, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd1, 5'd2, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd1, 5'd3, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd1, 5'd4, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd1, 5'd5, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd1, 5'd6, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd1, 5'd7, 1'd1} : pll_rate_sel_expected = 4'b0001;
  {PCIE, 4'd2, 5'd0, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd2, 5'd1, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd2, 5'd2, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd2, 5'd3, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd2, 5'd4, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd2, 5'd5, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd2, 5'd6, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd2, 5'd7, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd3, 5'd0, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd3, 5'd1, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd3, 5'd2, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd3, 5'd3, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd3, 5'd4, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd3, 5'd5, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd3, 5'd6, 1'd1} : pll_rate_sel_expected = 4'b0000;
  {PCIE, 4'd3, 5'd7, 1'd1} : pll_rate_sel_expected = 4'b0000;
default: pll_rate_sel_expected = 4'bzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel} )
  {USB, 4'd1, 5'd0, 1'd0} : fbdiv_expected = 10'b0110010000;
  {USB, 4'd1, 5'd1, 1'd0} : fbdiv_expected = 10'b0101001101;
  {USB, 4'd1, 5'd2, 1'd0} : fbdiv_expected = 10'b0011111010;
  {USB, 4'd1, 5'd3, 1'd0} : fbdiv_expected = 10'b0011001000;
  {USB, 4'd1, 5'd4, 1'd0} : fbdiv_expected = 10'b0010100000;
  {USB, 4'd1, 5'd5, 1'd0} : fbdiv_expected = 10'b0011001000;
  {USB, 4'd1, 5'd6, 1'd0} : fbdiv_expected = 10'b0001010000;
  {USB, 4'd1, 5'd7, 1'd0} : fbdiv_expected = 10'b0010000000;
  {USB, 4'd2, 5'd0, 1'd0} : fbdiv_expected = 10'b0110010000;
  {USB, 4'd2, 5'd1, 1'd0} : fbdiv_expected = 10'b0101001101;
  {USB, 4'd2, 5'd2, 1'd0} : fbdiv_expected = 10'b0011111010;
  {USB, 4'd2, 5'd3, 1'd0} : fbdiv_expected = 10'b0011001000;
  {USB, 4'd2, 5'd4, 1'd0} : fbdiv_expected = 10'b0010100000;
  {USB, 4'd2, 5'd5, 1'd0} : fbdiv_expected = 10'b0011001000;
  {USB, 4'd2, 5'd6, 1'd0} : fbdiv_expected = 10'b0001010000;
  {USB, 4'd2, 5'd7, 1'd0} : fbdiv_expected = 10'b0010000000;
  {SERDES, 4'd0, 5'd0, 1'd0} : fbdiv_expected = 10'b0110010000;
  {SERDES, 4'd0, 5'd1, 1'd0} : fbdiv_expected = 10'b0101001101;
  {SERDES, 4'd0, 5'd2, 1'd0} : fbdiv_expected = 10'b0011111010;
  {SERDES, 4'd0, 5'd3, 1'd0} : fbdiv_expected = 10'b0011001000;
  {SERDES, 4'd0, 5'd4, 1'd0} : fbdiv_expected = 10'b0010100000;
  {SERDES, 4'd0, 5'd5, 1'd0} : fbdiv_expected = 10'b0001100100;
  {SERDES, 4'd0, 5'd6, 1'd0} : fbdiv_expected = 10'b0001010000;
  {SERDES, 4'd0, 5'd7, 1'd0} : fbdiv_expected = 10'b0001000000;
  {SERDES, 4'd1, 5'd0, 1'd0} : fbdiv_expected = 10'b0111110100;
  {SERDES, 4'd1, 5'd1, 1'd0} : fbdiv_expected = 10'b0110100001;
  {SERDES, 4'd1, 5'd2, 1'd0} : fbdiv_expected = 10'b0100111001;
  {SERDES, 4'd1, 5'd3, 1'd0} : fbdiv_expected = 10'b0011111010;
  {SERDES, 4'd1, 5'd4, 1'd0} : fbdiv_expected = 10'b0011001000;
  {SERDES, 4'd1, 5'd5, 1'd0} : fbdiv_expected = 10'b0001111101;
  {SERDES, 4'd1, 5'd6, 1'd0} : fbdiv_expected = 10'b0001100100;
  {SERDES, 4'd1, 5'd7, 1'd0} : fbdiv_expected = 10'b0001010000;
  {SERDES, 4'd2, 5'd0, 1'd0} : fbdiv_expected = 10'b0110011101;
  {SERDES, 4'd2, 5'd1, 1'd0} : fbdiv_expected = 10'b0101011000;
  {SERDES, 4'd2, 5'd2, 1'd0} : fbdiv_expected = 10'b0100000010;
  {SERDES, 4'd2, 5'd3, 1'd0} : fbdiv_expected = 10'b0011001110;
  {SERDES, 4'd2, 5'd4, 1'd0} : fbdiv_expected = 10'b0010100101;
  {SERDES, 4'd2, 5'd5, 1'd0} : fbdiv_expected = 10'b0011001110;
  {SERDES, 4'd2, 5'd6, 1'd0} : fbdiv_expected = 10'b0010100101;
  {SERDES, 4'd2, 5'd7, 1'd0} : fbdiv_expected = 10'b0010000100;
  {SERDES, 4'd3, 5'd0, 1'd0} : fbdiv_expected = 10'b0111110100;
  {SERDES, 4'd3, 5'd1, 1'd0} : fbdiv_expected = 10'b0110100001;
  {SERDES, 4'd3, 5'd2, 1'd0} : fbdiv_expected = 10'b0100111001;
  {SERDES, 4'd3, 5'd3, 1'd0} : fbdiv_expected = 10'b0011111010;
  {SERDES, 4'd3, 5'd4, 1'd0} : fbdiv_expected = 10'b0011001000;
  {SERDES, 4'd3, 5'd5, 1'd0} : fbdiv_expected = 10'b0001111101;
  {SERDES, 4'd3, 5'd6, 1'd0} : fbdiv_expected = 10'b0001100100;
  {SERDES, 4'd3, 5'd7, 1'd0} : fbdiv_expected = 10'b0001010000;
  {SERDES, 4'd4, 5'd0, 1'd0} : fbdiv_expected = 10'b0110011101;
  {SERDES, 4'd4, 5'd1, 1'd0} : fbdiv_expected = 10'b0101011000;
  {SERDES, 4'd4, 5'd2, 1'd0} : fbdiv_expected = 10'b0100000010;
  {SERDES, 4'd4, 5'd3, 1'd0} : fbdiv_expected = 10'b0011001110;
  {SERDES, 4'd4, 5'd4, 1'd0} : fbdiv_expected = 10'b0010100101;
  {SERDES, 4'd4, 5'd5, 1'd0} : fbdiv_expected = 10'b0011001110;
  {SERDES, 4'd4, 5'd6, 1'd0} : fbdiv_expected = 10'b0010100101;
  {SERDES, 4'd4, 5'd7, 1'd0} : fbdiv_expected = 10'b0010000100;
  {SERDES, 4'd5, 5'd0, 1'd0} : fbdiv_expected = 10'b0111101000;
  {SERDES, 4'd5, 5'd1, 1'd0} : fbdiv_expected = 10'b0110010110;
  {SERDES, 4'd5, 5'd2, 1'd0} : fbdiv_expected = 10'b0100110001;
  {SERDES, 4'd5, 5'd3, 1'd0} : fbdiv_expected = 10'b0011110100;
  {SERDES, 4'd5, 5'd4, 1'd0} : fbdiv_expected = 10'b0011000011;
  {SERDES, 4'd5, 5'd5, 1'd0} : fbdiv_expected = 10'b0001111010;
  {SERDES, 4'd5, 5'd6, 1'd0} : fbdiv_expected = 10'b0011000011;
  {SERDES, 4'd5, 5'd7, 1'd0} : fbdiv_expected = 10'b0001001110;
  {SERDES, 4'd6, 5'd0, 1'd0} : fbdiv_expected = 10'b0111110100;
  {SERDES, 4'd6, 5'd1, 1'd0} : fbdiv_expected = 10'b0110100001;
  {SERDES, 4'd6, 5'd2, 1'd0} : fbdiv_expected = 10'b0100111001;
  {SERDES, 4'd6, 5'd3, 1'd0} : fbdiv_expected = 10'b0011111010;
  {SERDES, 4'd6, 5'd4, 1'd0} : fbdiv_expected = 10'b0011001000;
  {SERDES, 4'd6, 5'd5, 1'd0} : fbdiv_expected = 10'b0001111101;
  {SERDES, 4'd6, 5'd6, 1'd0} : fbdiv_expected = 10'b0001100100;
  {SERDES, 4'd6, 5'd7, 1'd0} : fbdiv_expected = 10'b0001010000;
  {SERDES, 4'd7, 5'd0, 1'd0} : fbdiv_expected = 10'b1000000100;
  {SERDES, 4'd7, 5'd1, 1'd0} : fbdiv_expected = 10'b0110101110;
  {SERDES, 4'd7, 5'd2, 1'd0} : fbdiv_expected = 10'b0101000010;
  {SERDES, 4'd7, 5'd3, 1'd0} : fbdiv_expected = 10'b0100000010;
  {SERDES, 4'd7, 5'd4, 1'd0} : fbdiv_expected = 10'b0011001110;
  {SERDES, 4'd7, 5'd5, 1'd0} : fbdiv_expected = 10'b0010000001;
  {SERDES, 4'd7, 5'd6, 1'd0} : fbdiv_expected = 10'b0001100111;
  {SERDES, 4'd7, 5'd7, 1'd0} : fbdiv_expected = 10'b0010100101;
  {SERDES, 4'd8, 5'd0, 1'd0} : fbdiv_expected = 10'b1000100110;
  {SERDES, 4'd8, 5'd1, 1'd0} : fbdiv_expected = 10'b0111001010;
  {SERDES, 4'd8, 5'd2, 1'd0} : fbdiv_expected = 10'b0101011000;
  {SERDES, 4'd8, 5'd3, 1'd0} : fbdiv_expected = 10'b0100010011;
  {SERDES, 4'd8, 5'd4, 1'd0} : fbdiv_expected = 10'b0011011100;
  {SERDES, 4'd8, 5'd5, 1'd0} : fbdiv_expected = 10'b0100010011;
  {SERDES, 4'd8, 5'd6, 1'd0} : fbdiv_expected = 10'b0011011100;
  {SERDES, 4'd8, 5'd7, 1'd0} : fbdiv_expected = 10'b0010110000;
  {SERDES, 4'd9, 5'd0, 1'd0} : fbdiv_expected = 10'b1000110011;
  {SERDES, 4'd9, 5'd1, 1'd0} : fbdiv_expected = 10'b0111010101;
  {SERDES, 4'd9, 5'd2, 1'd0} : fbdiv_expected = 10'b0101100000;
  {SERDES, 4'd9, 5'd3, 1'd0} : fbdiv_expected = 10'b0100011001;
  {SERDES, 4'd9, 5'd4, 1'd0} : fbdiv_expected = 10'b0011100001;
  {SERDES, 4'd9, 5'd5, 1'd0} : fbdiv_expected = 10'b0100011001;
  {SERDES, 4'd9, 5'd6, 1'd0} : fbdiv_expected = 10'b0011100001;
  {SERDES, 4'd9, 5'd7, 1'd0} : fbdiv_expected = 10'b0010110100;
  {SERDES, 4'd12, 5'd0, 1'd0} : fbdiv_expected = 10'b0110010000;
  {SERDES, 4'd12, 5'd1, 1'd0} : fbdiv_expected = 10'b0101001101;
  {SERDES, 4'd12, 5'd2, 1'd0} : fbdiv_expected = 10'b0011111010;
  {SERDES, 4'd12, 5'd3, 1'd0} : fbdiv_expected = 10'b0011001000;
  {SERDES, 4'd12, 5'd4, 1'd0} : fbdiv_expected = 10'b0010100000;
  {SERDES, 4'd12, 5'd5, 1'd0} : fbdiv_expected = 10'b0001100100;
  {SERDES, 4'd12, 5'd6, 1'd0} : fbdiv_expected = 10'b0001010000;
  {SERDES, 4'd12, 5'd7, 1'd0} : fbdiv_expected = 10'b0001000000;
  {SERDES, 4'd13, 5'd0, 1'd0} : fbdiv_expected = 10'b0110011101;
  {SERDES, 4'd13, 5'd1, 1'd0} : fbdiv_expected = 10'b0101011000;
  {SERDES, 4'd13, 5'd2, 1'd0} : fbdiv_expected = 10'b0100000010;
  {SERDES, 4'd13, 5'd3, 1'd0} : fbdiv_expected = 10'b0011001110;
  {SERDES, 4'd13, 5'd4, 1'd0} : fbdiv_expected = 10'b0010100101;
  {SERDES, 4'd13, 5'd5, 1'd0} : fbdiv_expected = 10'b0011001110;
  {SERDES, 4'd13, 5'd6, 1'd0} : fbdiv_expected = 10'b0010100101;
  {SERDES, 4'd13, 5'd7, 1'd0} : fbdiv_expected = 10'b0010000100;
  {SAS, 4'd0, 5'd0, 1'd0} : fbdiv_expected = 10'b0111100000;
  {SAS, 4'd0, 5'd1, 1'd0} : fbdiv_expected = 10'b0110010000;
  {SAS, 4'd0, 5'd2, 1'd0} : fbdiv_expected = 10'b0100101100;
  {SAS, 4'd0, 5'd3, 1'd0} : fbdiv_expected = 10'b0011110000;
  {SAS, 4'd0, 5'd4, 1'd0} : fbdiv_expected = 10'b0011000000;
  {SAS, 4'd0, 5'd5, 1'd0} : fbdiv_expected = 10'b0011110000;
  {SAS, 4'd0, 5'd6, 1'd0} : fbdiv_expected = 10'b0001100000;
  {SAS, 4'd0, 5'd7, 1'd0} : fbdiv_expected = 10'b0100110011;
  {SAS, 4'd1, 5'd0, 1'd0} : fbdiv_expected = 10'b0111100000;
  {SAS, 4'd1, 5'd1, 1'd0} : fbdiv_expected = 10'b0110010000;
  {SAS, 4'd1, 5'd2, 1'd0} : fbdiv_expected = 10'b0100101100;
  {SAS, 4'd1, 5'd3, 1'd0} : fbdiv_expected = 10'b0011110000;
  {SAS, 4'd1, 5'd4, 1'd0} : fbdiv_expected = 10'b0011000000;
  {SAS, 4'd1, 5'd5, 1'd0} : fbdiv_expected = 10'b0011110000;
  {SAS, 4'd1, 5'd6, 1'd0} : fbdiv_expected = 10'b0001100000;
  {SAS, 4'd1, 5'd7, 1'd0} : fbdiv_expected = 10'b0100110011;
  {SAS, 4'd2, 5'd0, 1'd0} : fbdiv_expected = 10'b0111100000;
  {SAS, 4'd2, 5'd1, 1'd0} : fbdiv_expected = 10'b0110010000;
  {SAS, 4'd2, 5'd2, 1'd0} : fbdiv_expected = 10'b0100101100;
  {SAS, 4'd2, 5'd3, 1'd0} : fbdiv_expected = 10'b0011110000;
  {SAS, 4'd2, 5'd4, 1'd0} : fbdiv_expected = 10'b0011000000;
  {SAS, 4'd2, 5'd5, 1'd0} : fbdiv_expected = 10'b0011110000;
  {SAS, 4'd2, 5'd6, 1'd0} : fbdiv_expected = 10'b0001100000;
  {SAS, 4'd2, 5'd7, 1'd0} : fbdiv_expected = 10'b0100110011;
  {SAS, 4'd3, 5'd0, 1'd0} : fbdiv_expected = 10'b0111100000;
  {SAS, 4'd3, 5'd1, 1'd0} : fbdiv_expected = 10'b0110010000;
  {SAS, 4'd3, 5'd2, 1'd0} : fbdiv_expected = 10'b0100101100;
  {SAS, 4'd3, 5'd3, 1'd0} : fbdiv_expected = 10'b0011110000;
  {SAS, 4'd3, 5'd4, 1'd0} : fbdiv_expected = 10'b0011000000;
  {SAS, 4'd3, 5'd5, 1'd0} : fbdiv_expected = 10'b0011110000;
  {SAS, 4'd3, 5'd6, 1'd0} : fbdiv_expected = 10'b0001100000;
  {SAS, 4'd3, 5'd7, 1'd0} : fbdiv_expected = 10'b0100110011;
  {SAS, 4'd4, 5'd0, 1'd0} : fbdiv_expected = 10'b0111000010;
  {SAS, 4'd4, 5'd1, 1'd0} : fbdiv_expected = 10'b0101110111;
  {SAS, 4'd4, 5'd2, 1'd0} : fbdiv_expected = 10'b0100011001;
  {SAS, 4'd4, 5'd3, 1'd0} : fbdiv_expected = 10'b0011100001;
  {SAS, 4'd4, 5'd4, 1'd0} : fbdiv_expected = 10'b0101101000;
  {SAS, 4'd4, 5'd5, 1'd0} : fbdiv_expected = 10'b0011100001;
  {SAS, 4'd4, 5'd6, 1'd0} : fbdiv_expected = 10'b0001011010;
  {SAS, 4'd4, 5'd7, 1'd0} : fbdiv_expected = 10'b0010010000;
  {PCIE, 4'd2, 5'd0, 1'd0} : fbdiv_expected = 10'b0101000000;
  {PCIE, 4'd2, 5'd1, 1'd0} : fbdiv_expected = 10'b0100001011;
  {PCIE, 4'd2, 5'd2, 1'd0} : fbdiv_expected = 10'b0011001000;
  {PCIE, 4'd2, 5'd3, 1'd0} : fbdiv_expected = 10'b0101000000;
  {PCIE, 4'd2, 5'd4, 1'd0} : fbdiv_expected = 10'b0010000000;
  {PCIE, 4'd2, 5'd5, 1'd0} : fbdiv_expected = 10'b0001010000;
  {PCIE, 4'd2, 5'd6, 1'd0} : fbdiv_expected = 10'b0001000000;
  {PCIE, 4'd2, 5'd7, 1'd0} : fbdiv_expected = 10'b0011001101;
  {PCIE, 4'd3, 5'd0, 1'd0} : fbdiv_expected = 10'b0101000000;
  {PCIE, 4'd3, 5'd1, 1'd0} : fbdiv_expected = 10'b0100001011;
  {PCIE, 4'd3, 5'd2, 1'd0} : fbdiv_expected = 10'b0011001000;
  {PCIE, 4'd3, 5'd3, 1'd0} : fbdiv_expected = 10'b0101000000;
  {PCIE, 4'd3, 5'd4, 1'd0} : fbdiv_expected = 10'b0010000000;
  {PCIE, 4'd3, 5'd5, 1'd0} : fbdiv_expected = 10'b0001010000;
  {PCIE, 4'd3, 5'd6, 1'd0} : fbdiv_expected = 10'b0001000000;
  {PCIE, 4'd3, 5'd7, 1'd0} : fbdiv_expected = 10'b0011001101;
  {USB, 4'd1, 5'd0, 1'd1} : fbdiv_expected = 10'b0001100100;
  {USB, 4'd1, 5'd1, 1'd1} : fbdiv_expected = 10'b0001010011;
  {USB, 4'd1, 5'd2, 1'd1} : fbdiv_expected = 10'b0001111101;
  {USB, 4'd1, 5'd3, 1'd1} : fbdiv_expected = 10'b0000110010;
  {USB, 4'd1, 5'd4, 1'd1} : fbdiv_expected = 10'b0000101000;
  {USB, 4'd1, 5'd5, 1'd1} : fbdiv_expected = 10'b0000110010;
  {USB, 4'd1, 5'd6, 1'd1} : fbdiv_expected = 10'b0000010100;
  {USB, 4'd1, 5'd7, 1'd1} : fbdiv_expected = 10'b0000100000;
  {USB, 4'd2, 5'd0, 1'd1} : fbdiv_expected = 10'b0001100100;
  {USB, 4'd2, 5'd1, 1'd1} : fbdiv_expected = 10'b0001010011;
  {USB, 4'd2, 5'd2, 1'd1} : fbdiv_expected = 10'b0001111101;
  {USB, 4'd2, 5'd3, 1'd1} : fbdiv_expected = 10'b0000110010;
  {USB, 4'd2, 5'd4, 1'd1} : fbdiv_expected = 10'b0000101000;
  {USB, 4'd2, 5'd5, 1'd1} : fbdiv_expected = 10'b0000110010;
  {USB, 4'd2, 5'd6, 1'd1} : fbdiv_expected = 10'b0000010100;
  {USB, 4'd2, 5'd7, 1'd1} : fbdiv_expected = 10'b0000100000;
  {SERDES, 4'd0, 5'd0, 1'd1} : fbdiv_expected = 10'b0001100100;
  {SERDES, 4'd0, 5'd1, 1'd1} : fbdiv_expected = 10'b0001010011;
  {SERDES, 4'd0, 5'd2, 1'd1} : fbdiv_expected = 10'b0001111101;
  {SERDES, 4'd0, 5'd3, 1'd1} : fbdiv_expected = 10'b0001100100;
  {SERDES, 4'd0, 5'd4, 1'd1} : fbdiv_expected = 10'b0001111000;
  {SERDES, 4'd0, 5'd5, 1'd1} : fbdiv_expected = 10'b0001001011;
  {SERDES, 4'd0, 5'd6, 1'd1} : fbdiv_expected = 10'b0000111100;
  {SERDES, 4'd0, 5'd7, 1'd1} : fbdiv_expected = 10'b0000100000;
  {SERDES, 4'd1, 5'd0, 1'd1} : fbdiv_expected = 10'b0001111101;
  {SERDES, 4'd1, 5'd1, 1'd1} : fbdiv_expected = 10'b0001101000;
  {SERDES, 4'd1, 5'd2, 1'd1} : fbdiv_expected = 10'b0001001110;
  {SERDES, 4'd1, 5'd3, 1'd1} : fbdiv_expected = 10'b0001111101;
  {SERDES, 4'd1, 5'd4, 1'd1} : fbdiv_expected = 10'b0000110010;
  {SERDES, 4'd1, 5'd5, 1'd1} : fbdiv_expected = 10'b0001011110;
  {SERDES, 4'd1, 5'd6, 1'd1} : fbdiv_expected = 10'b0000011001;
  {SERDES, 4'd1, 5'd7, 1'd1} : fbdiv_expected = 10'b0000010100;
  {SERDES, 4'd2, 5'd0, 1'd1} : fbdiv_expected = 10'b0001100111;
  {SERDES, 4'd2, 5'd1, 1'd1} : fbdiv_expected = 10'b0010101100;
  {SERDES, 4'd2, 5'd2, 1'd1} : fbdiv_expected = 10'b0011000001;
  {SERDES, 4'd2, 5'd3, 1'd1} : fbdiv_expected = 10'b0001100111;
  {SERDES, 4'd2, 5'd4, 1'd1} : fbdiv_expected = 10'b0010100101;
  {SERDES, 4'd2, 5'd5, 1'd1} : fbdiv_expected = 10'b0001100111;
  {SERDES, 4'd2, 5'd6, 1'd1} : fbdiv_expected = 10'b0000111110;
  {SERDES, 4'd2, 5'd7, 1'd1} : fbdiv_expected = 10'b0000100001;
  {SERDES, 4'd3, 5'd0, 1'd1} : fbdiv_expected = 10'b0001111101;
  {SERDES, 4'd3, 5'd1, 1'd1} : fbdiv_expected = 10'b0001101000;
  {SERDES, 4'd3, 5'd2, 1'd1} : fbdiv_expected = 10'b0001001110;
  {SERDES, 4'd3, 5'd3, 1'd1} : fbdiv_expected = 10'b0001111101;
  {SERDES, 4'd3, 5'd4, 1'd1} : fbdiv_expected = 10'b0000110010;
  {SERDES, 4'd3, 5'd5, 1'd1} : fbdiv_expected = 10'b0001011110;
  {SERDES, 4'd3, 5'd6, 1'd1} : fbdiv_expected = 10'b0000011001;
  {SERDES, 4'd3, 5'd7, 1'd1} : fbdiv_expected = 10'b0000010100;
  {SERDES, 4'd4, 5'd0, 1'd1} : fbdiv_expected = 10'b0001100111;
  {SERDES, 4'd4, 5'd1, 1'd1} : fbdiv_expected = 10'b0010101100;
  {SERDES, 4'd4, 5'd2, 1'd1} : fbdiv_expected = 10'b0011000001;
  {SERDES, 4'd4, 5'd3, 1'd1} : fbdiv_expected = 10'b0001100111;
  {SERDES, 4'd4, 5'd4, 1'd1} : fbdiv_expected = 10'b0010100101;
  {SERDES, 4'd4, 5'd5, 1'd1} : fbdiv_expected = 10'b0001100111;
  {SERDES, 4'd4, 5'd6, 1'd1} : fbdiv_expected = 10'b0000111110;
  {SERDES, 4'd4, 5'd7, 1'd1} : fbdiv_expected = 10'b0000100001;
  {SERDES, 4'd5, 5'd0, 1'd1} : fbdiv_expected = 10'b0001111010;
  {SERDES, 4'd5, 5'd1, 1'd1} : fbdiv_expected = 10'b0011001011;
  {SERDES, 4'd5, 5'd2, 1'd1} : fbdiv_expected = 10'b0001001100;
  {SERDES, 4'd5, 5'd3, 1'd1} : fbdiv_expected = 10'b0001111010;
  {SERDES, 4'd5, 5'd4, 1'd1} : fbdiv_expected = 10'b0000110001;
  {SERDES, 4'd5, 5'd5, 1'd1} : fbdiv_expected = 10'b0000111101;
  {SERDES, 4'd5, 5'd6, 1'd1} : fbdiv_expected = 10'b0000110001;
  {SERDES, 4'd5, 5'd7, 1'd1} : fbdiv_expected = 10'b0000100111;
  {SERDES, 4'd6, 5'd0, 1'd1} : fbdiv_expected = 10'b0001111101;
  {SERDES, 4'd6, 5'd1, 1'd1} : fbdiv_expected = 10'b0001101000;
  {SERDES, 4'd6, 5'd2, 1'd1} : fbdiv_expected = 10'b0001001110;
  {SERDES, 4'd6, 5'd3, 1'd1} : fbdiv_expected = 10'b0001111101;
  {SERDES, 4'd6, 5'd4, 1'd1} : fbdiv_expected = 10'b0000110010;
  {SERDES, 4'd6, 5'd5, 1'd1} : fbdiv_expected = 10'b0001011110;
  {SERDES, 4'd6, 5'd6, 1'd1} : fbdiv_expected = 10'b0000011001;
  {SERDES, 4'd6, 5'd7, 1'd1} : fbdiv_expected = 10'b0000010100;
  {SERDES, 4'd7, 5'd0, 1'd1} : fbdiv_expected = 10'b0010000001;
  {SERDES, 4'd7, 5'd1, 1'd1} : fbdiv_expected = 10'b0001101011;
  {SERDES, 4'd7, 5'd2, 1'd1} : fbdiv_expected = 10'b0001010001;
  {SERDES, 4'd7, 5'd3, 1'd1} : fbdiv_expected = 10'b0010000001;
  {SERDES, 4'd7, 5'd4, 1'd1} : fbdiv_expected = 10'b0010011011;
  {SERDES, 4'd7, 5'd5, 1'd1} : fbdiv_expected = 10'b0001100001;
  {SERDES, 4'd7, 5'd6, 1'd1} : fbdiv_expected = 10'b0010000001;
  {SERDES, 4'd7, 5'd7, 1'd1} : fbdiv_expected = 10'b0000111110;
  {SERDES, 4'd8, 5'd0, 1'd1} : fbdiv_expected = 10'b0010001010;
  {SERDES, 4'd8, 5'd1, 1'd1} : fbdiv_expected = 10'b0011100101;
  {SERDES, 4'd8, 5'd2, 1'd1} : fbdiv_expected = 10'b0001010110;
  {SERDES, 4'd8, 5'd3, 1'd1} : fbdiv_expected = 10'b0001000101;
  {SERDES, 4'd8, 5'd4, 1'd1} : fbdiv_expected = 10'b0000110111;
  {SERDES, 4'd8, 5'd5, 1'd1} : fbdiv_expected = 10'b0001000101;
  {SERDES, 4'd8, 5'd6, 1'd1} : fbdiv_expected = 10'b0000110111;
  {SERDES, 4'd8, 5'd7, 1'd1} : fbdiv_expected = 10'b0000101100;
  {SERDES, 4'd9, 5'd0, 1'd1} : fbdiv_expected = 10'b0010001101;
  {SERDES, 4'd9, 5'd1, 1'd1} : fbdiv_expected = 10'b0001110101;
  {SERDES, 4'd9, 5'd2, 1'd1} : fbdiv_expected = 10'b0001011000;
  {SERDES, 4'd9, 5'd3, 1'd1} : fbdiv_expected = 10'b0001000110;
  {SERDES, 4'd9, 5'd4, 1'd1} : fbdiv_expected = 10'b0000111000;
  {SERDES, 4'd9, 5'd5, 1'd1} : fbdiv_expected = 10'b0001000110;
  {SERDES, 4'd9, 5'd6, 1'd1} : fbdiv_expected = 10'b0000111000;
  {SERDES, 4'd9, 5'd7, 1'd1} : fbdiv_expected = 10'b0000101101;
  {SERDES, 4'd12, 5'd0, 1'd1} : fbdiv_expected = 10'b0001100100;
  {SERDES, 4'd12, 5'd1, 1'd1} : fbdiv_expected = 10'b0001010011;
  {SERDES, 4'd12, 5'd2, 1'd1} : fbdiv_expected = 10'b0001111101;
  {SERDES, 4'd12, 5'd3, 1'd1} : fbdiv_expected = 10'b0001100100;
  {SERDES, 4'd12, 5'd4, 1'd1} : fbdiv_expected = 10'b0001111000;
  {SERDES, 4'd12, 5'd5, 1'd1} : fbdiv_expected = 10'b0001001011;
  {SERDES, 4'd12, 5'd6, 1'd1} : fbdiv_expected = 10'b0000111100;
  {SERDES, 4'd12, 5'd7, 1'd1} : fbdiv_expected = 10'b0000100000;
  {SERDES, 4'd13, 5'd0, 1'd1} : fbdiv_expected = 10'b0001100111;
  {SERDES, 4'd13, 5'd1, 1'd1} : fbdiv_expected = 10'b0010101100;
  {SERDES, 4'd13, 5'd2, 1'd1} : fbdiv_expected = 10'b0011000001;
  {SERDES, 4'd13, 5'd3, 1'd1} : fbdiv_expected = 10'b0001100111;
  {SERDES, 4'd13, 5'd4, 1'd1} : fbdiv_expected = 10'b0010100101;
  {SERDES, 4'd13, 5'd5, 1'd1} : fbdiv_expected = 10'b0001100111;
  {SERDES, 4'd13, 5'd6, 1'd1} : fbdiv_expected = 10'b0000111110;
  {SERDES, 4'd13, 5'd7, 1'd1} : fbdiv_expected = 10'b0000100001;
  {SAS, 4'd0, 5'd0, 1'd1} : fbdiv_expected = 10'b0001111000;
  {SAS, 4'd0, 5'd1, 1'd1} : fbdiv_expected = 10'b0001100100;
  {SAS, 4'd0, 5'd2, 1'd1} : fbdiv_expected = 10'b0011100010;
  {SAS, 4'd0, 5'd3, 1'd1} : fbdiv_expected = 10'b0010110101;
  {SAS, 4'd0, 5'd4, 1'd1} : fbdiv_expected = 10'b0000110000;
  {SAS, 4'd0, 5'd5, 1'd1} : fbdiv_expected = 10'b0000111100;
  {SAS, 4'd0, 5'd6, 1'd1} : fbdiv_expected = 10'b0000011000;
  {SAS, 4'd0, 5'd7, 1'd1} : fbdiv_expected = 10'b0001001101;
  {SAS, 4'd1, 5'd0, 1'd1} : fbdiv_expected = 10'b0001111000;
  {SAS, 4'd1, 5'd1, 1'd1} : fbdiv_expected = 10'b0001100100;
  {SAS, 4'd1, 5'd2, 1'd1} : fbdiv_expected = 10'b0011100010;
  {SAS, 4'd1, 5'd3, 1'd1} : fbdiv_expected = 10'b0010110101;
  {SAS, 4'd1, 5'd4, 1'd1} : fbdiv_expected = 10'b0000110000;
  {SAS, 4'd1, 5'd5, 1'd1} : fbdiv_expected = 10'b0000111100;
  {SAS, 4'd1, 5'd6, 1'd1} : fbdiv_expected = 10'b0000011000;
  {SAS, 4'd1, 5'd7, 1'd1} : fbdiv_expected = 10'b0001001101;
  {SAS, 4'd2, 5'd0, 1'd1} : fbdiv_expected = 10'b0001111000;
  {SAS, 4'd2, 5'd1, 1'd1} : fbdiv_expected = 10'b0001100100;
  {SAS, 4'd2, 5'd2, 1'd1} : fbdiv_expected = 10'b0011100010;
  {SAS, 4'd2, 5'd3, 1'd1} : fbdiv_expected = 10'b0010110101;
  {SAS, 4'd2, 5'd4, 1'd1} : fbdiv_expected = 10'b0000110000;
  {SAS, 4'd2, 5'd5, 1'd1} : fbdiv_expected = 10'b0000111100;
  {SAS, 4'd2, 5'd6, 1'd1} : fbdiv_expected = 10'b0000011000;
  {SAS, 4'd2, 5'd7, 1'd1} : fbdiv_expected = 10'b0001001101;
  {SAS, 4'd3, 5'd0, 1'd1} : fbdiv_expected = 10'b0001111000;
  {SAS, 4'd3, 5'd1, 1'd1} : fbdiv_expected = 10'b0001100100;
  {SAS, 4'd3, 5'd2, 1'd1} : fbdiv_expected = 10'b0011100010;
  {SAS, 4'd3, 5'd3, 1'd1} : fbdiv_expected = 10'b0010110101;
  {SAS, 4'd3, 5'd4, 1'd1} : fbdiv_expected = 10'b0000110000;
  {SAS, 4'd3, 5'd5, 1'd1} : fbdiv_expected = 10'b0000111100;
  {SAS, 4'd3, 5'd6, 1'd1} : fbdiv_expected = 10'b0000011000;
  {SAS, 4'd3, 5'd7, 1'd1} : fbdiv_expected = 10'b0001001101;
  {SAS, 4'd4, 5'd0, 1'd1} : fbdiv_expected = 10'b0001110001;
  {SAS, 4'd4, 5'd1, 1'd1} : fbdiv_expected = 10'b0001011110;
  {SAS, 4'd4, 5'd2, 1'd1} : fbdiv_expected = 10'b0001000110;
  {SAS, 4'd4, 5'd3, 1'd1} : fbdiv_expected = 10'b0000111000;
  {SAS, 4'd4, 5'd4, 1'd1} : fbdiv_expected = 10'b0001011010;
  {SAS, 4'd4, 5'd5, 1'd1} : fbdiv_expected = 10'b0000111000;
  {SAS, 4'd4, 5'd6, 1'd1} : fbdiv_expected = 10'b0000101101;
  {SAS, 4'd4, 5'd7, 1'd1} : fbdiv_expected = 10'b0000100100;
  {PCIE, 4'd2, 5'd0, 1'd1} : fbdiv_expected = 10'b0001010000;
  {PCIE, 4'd2, 5'd1, 1'd1} : fbdiv_expected = 10'b0010000101;
  {PCIE, 4'd2, 5'd2, 1'd1} : fbdiv_expected = 10'b0000110010;
  {PCIE, 4'd2, 5'd3, 1'd1} : fbdiv_expected = 10'b0001010000;
  {PCIE, 4'd2, 5'd4, 1'd1} : fbdiv_expected = 10'b0000100000;
  {PCIE, 4'd2, 5'd5, 1'd1} : fbdiv_expected = 10'b0000010100;
  {PCIE, 4'd2, 5'd6, 1'd1} : fbdiv_expected = 10'b0000010000;
  {PCIE, 4'd2, 5'd7, 1'd1} : fbdiv_expected = 10'b0000110011;
  {PCIE, 4'd3, 5'd0, 1'd1} : fbdiv_expected = 10'b0001010000;
  {PCIE, 4'd3, 5'd1, 1'd1} : fbdiv_expected = 10'b0010000101;
  {PCIE, 4'd3, 5'd2, 1'd1} : fbdiv_expected = 10'b0000110010;
  {PCIE, 4'd3, 5'd3, 1'd1} : fbdiv_expected = 10'b0001010000;
  {PCIE, 4'd3, 5'd4, 1'd1} : fbdiv_expected = 10'b0000100000;
  {PCIE, 4'd3, 5'd5, 1'd1} : fbdiv_expected = 10'b0000010100;
  {PCIE, 4'd3, 5'd6, 1'd1} : fbdiv_expected = 10'b0000010000;
  {PCIE, 4'd3, 5'd7, 1'd1} : fbdiv_expected = 10'b0000110011;
default: fbdiv_expected = 10'bzzzzzzzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel} )
  {USB, 4'd1, 5'd0, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd1, 5'd1, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd1, 5'd2, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd1, 5'd3, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd1, 5'd4, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd1, 5'd5, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd1, 5'd6, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd1, 5'd7, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd2, 5'd0, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd2, 5'd1, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd2, 5'd2, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd2, 5'd3, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd2, 5'd4, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd2, 5'd5, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd2, 5'd6, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd2, 5'd7, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd0, 5'd0, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd0, 5'd1, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd0, 5'd2, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd0, 5'd3, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd0, 5'd4, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd0, 5'd5, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd0, 5'd6, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd0, 5'd7, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd1, 5'd0, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd1, 5'd1, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd1, 5'd2, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd1, 5'd3, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd1, 5'd4, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd1, 5'd5, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd1, 5'd6, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd1, 5'd7, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd2, 5'd0, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd2, 5'd1, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd2, 5'd2, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd2, 5'd3, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd2, 5'd4, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd2, 5'd5, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd2, 5'd6, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd2, 5'd7, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd3, 5'd0, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd3, 5'd1, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd3, 5'd2, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd3, 5'd3, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd3, 5'd4, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd3, 5'd5, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd3, 5'd6, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd3, 5'd7, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd4, 5'd0, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd4, 5'd1, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd4, 5'd2, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd4, 5'd3, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd4, 5'd4, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd4, 5'd5, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd4, 5'd6, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd4, 5'd7, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd5, 5'd0, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SERDES, 4'd5, 5'd1, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SERDES, 4'd5, 5'd2, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SERDES, 4'd5, 5'd3, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SERDES, 4'd5, 5'd4, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SERDES, 4'd5, 5'd5, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SERDES, 4'd5, 5'd6, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SERDES, 4'd5, 5'd7, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SERDES, 4'd6, 5'd0, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd6, 5'd1, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd6, 5'd2, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd6, 5'd3, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd6, 5'd4, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd6, 5'd5, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd6, 5'd6, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd6, 5'd7, 1'd0} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd7, 5'd0, 1'd0} : fbdiv_cal_expected = 10'b0000011010;
  {SERDES, 4'd7, 5'd1, 1'd0} : fbdiv_cal_expected = 10'b0000011010;
  {SERDES, 4'd7, 5'd2, 1'd0} : fbdiv_cal_expected = 10'b0000011010;
  {SERDES, 4'd7, 5'd3, 1'd0} : fbdiv_cal_expected = 10'b0000011010;
  {SERDES, 4'd7, 5'd4, 1'd0} : fbdiv_cal_expected = 10'b0000011010;
  {SERDES, 4'd7, 5'd5, 1'd0} : fbdiv_cal_expected = 10'b0000011010;
  {SERDES, 4'd7, 5'd6, 1'd0} : fbdiv_cal_expected = 10'b0000011010;
  {SERDES, 4'd7, 5'd7, 1'd0} : fbdiv_cal_expected = 10'b0000011010;
  {SERDES, 4'd8, 5'd0, 1'd0} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd8, 5'd1, 1'd0} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd8, 5'd2, 1'd0} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd8, 5'd3, 1'd0} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd8, 5'd4, 1'd0} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd8, 5'd5, 1'd0} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd8, 5'd6, 1'd0} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd8, 5'd7, 1'd0} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd9, 5'd0, 1'd0} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd9, 5'd1, 1'd0} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd9, 5'd2, 1'd0} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd9, 5'd3, 1'd0} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd9, 5'd4, 1'd0} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd9, 5'd5, 1'd0} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd9, 5'd6, 1'd0} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd9, 5'd7, 1'd0} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd12, 5'd0, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd12, 5'd1, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd12, 5'd2, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd12, 5'd3, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd12, 5'd4, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd12, 5'd5, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd12, 5'd6, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd12, 5'd7, 1'd0} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd13, 5'd0, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd13, 5'd1, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd13, 5'd2, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd13, 5'd3, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd13, 5'd4, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd13, 5'd5, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd13, 5'd6, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd13, 5'd7, 1'd0} : fbdiv_cal_expected = 10'b0000010101;
  {SAS, 4'd0, 5'd0, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd0, 5'd1, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd0, 5'd2, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd0, 5'd3, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd0, 5'd4, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd0, 5'd5, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd0, 5'd6, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd0, 5'd7, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd1, 5'd0, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd1, 5'd1, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd1, 5'd2, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd1, 5'd3, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd1, 5'd4, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd1, 5'd5, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd1, 5'd6, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd1, 5'd7, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd2, 5'd0, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd2, 5'd1, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd2, 5'd2, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd2, 5'd3, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd2, 5'd4, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd2, 5'd5, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd2, 5'd6, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd2, 5'd7, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd3, 5'd0, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd3, 5'd1, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd3, 5'd2, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd3, 5'd3, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd3, 5'd4, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd3, 5'd5, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd3, 5'd6, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd3, 5'd7, 1'd0} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd4, 5'd0, 1'd0} : fbdiv_cal_expected = 10'b0000010111;
  {SAS, 4'd4, 5'd1, 1'd0} : fbdiv_cal_expected = 10'b0000010111;
  {SAS, 4'd4, 5'd2, 1'd0} : fbdiv_cal_expected = 10'b0000010111;
  {SAS, 4'd4, 5'd3, 1'd0} : fbdiv_cal_expected = 10'b0000010111;
  {SAS, 4'd4, 5'd4, 1'd0} : fbdiv_cal_expected = 10'b0000010111;
  {SAS, 4'd4, 5'd5, 1'd0} : fbdiv_cal_expected = 10'b0000010111;
  {SAS, 4'd4, 5'd6, 1'd0} : fbdiv_cal_expected = 10'b0000010111;
  {SAS, 4'd4, 5'd7, 1'd0} : fbdiv_cal_expected = 10'b0000010111;
  {PCIE, 4'd2, 5'd0, 1'd0} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd2, 5'd1, 1'd0} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd2, 5'd2, 1'd0} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd2, 5'd3, 1'd0} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd2, 5'd4, 1'd0} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd2, 5'd5, 1'd0} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd2, 5'd6, 1'd0} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd2, 5'd7, 1'd0} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd3, 5'd0, 1'd0} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd3, 5'd1, 1'd0} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd3, 5'd2, 1'd0} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd3, 5'd3, 1'd0} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd3, 5'd4, 1'd0} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd3, 5'd5, 1'd0} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd3, 5'd6, 1'd0} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd3, 5'd7, 1'd0} : fbdiv_cal_expected = 10'b0000010000;
  {USB, 4'd1, 5'd0, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd1, 5'd1, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd1, 5'd2, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd1, 5'd3, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd1, 5'd4, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd1, 5'd5, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd1, 5'd6, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd1, 5'd7, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd2, 5'd0, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd2, 5'd1, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd2, 5'd2, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd2, 5'd3, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd2, 5'd4, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd2, 5'd5, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd2, 5'd6, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {USB, 4'd2, 5'd7, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd0, 5'd0, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd0, 5'd1, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd0, 5'd2, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd0, 5'd3, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd0, 5'd4, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd0, 5'd5, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd0, 5'd6, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd0, 5'd7, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd1, 5'd0, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd1, 5'd1, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd1, 5'd2, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd1, 5'd3, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd1, 5'd4, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd1, 5'd5, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd1, 5'd6, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd1, 5'd7, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd2, 5'd0, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd2, 5'd1, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd2, 5'd2, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd2, 5'd3, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd2, 5'd4, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd2, 5'd5, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd2, 5'd6, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd2, 5'd7, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd3, 5'd0, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd3, 5'd1, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd3, 5'd2, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd3, 5'd3, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd3, 5'd4, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd3, 5'd5, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd3, 5'd6, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd3, 5'd7, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd4, 5'd0, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd4, 5'd1, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd4, 5'd2, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd4, 5'd3, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd4, 5'd4, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd4, 5'd5, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd4, 5'd6, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd4, 5'd7, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd5, 5'd0, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SERDES, 4'd5, 5'd1, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SERDES, 4'd5, 5'd2, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SERDES, 4'd5, 5'd3, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SERDES, 4'd5, 5'd4, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SERDES, 4'd5, 5'd5, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SERDES, 4'd5, 5'd6, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SERDES, 4'd5, 5'd7, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SERDES, 4'd6, 5'd0, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd6, 5'd1, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd6, 5'd2, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd6, 5'd3, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd6, 5'd4, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd6, 5'd5, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd6, 5'd6, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd6, 5'd7, 1'd1} : fbdiv_cal_expected = 10'b0000011001;
  {SERDES, 4'd7, 5'd0, 1'd1} : fbdiv_cal_expected = 10'b0000011010;
  {SERDES, 4'd7, 5'd1, 1'd1} : fbdiv_cal_expected = 10'b0000011010;
  {SERDES, 4'd7, 5'd2, 1'd1} : fbdiv_cal_expected = 10'b0000011010;
  {SERDES, 4'd7, 5'd3, 1'd1} : fbdiv_cal_expected = 10'b0000011010;
  {SERDES, 4'd7, 5'd4, 1'd1} : fbdiv_cal_expected = 10'b0000011010;
  {SERDES, 4'd7, 5'd5, 1'd1} : fbdiv_cal_expected = 10'b0000011010;
  {SERDES, 4'd7, 5'd6, 1'd1} : fbdiv_cal_expected = 10'b0000011010;
  {SERDES, 4'd7, 5'd7, 1'd1} : fbdiv_cal_expected = 10'b0000011010;
  {SERDES, 4'd8, 5'd0, 1'd1} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd8, 5'd1, 1'd1} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd8, 5'd2, 1'd1} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd8, 5'd3, 1'd1} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd8, 5'd4, 1'd1} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd8, 5'd5, 1'd1} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd8, 5'd6, 1'd1} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd8, 5'd7, 1'd1} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd9, 5'd0, 1'd1} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd9, 5'd1, 1'd1} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd9, 5'd2, 1'd1} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd9, 5'd3, 1'd1} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd9, 5'd4, 1'd1} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd9, 5'd5, 1'd1} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd9, 5'd6, 1'd1} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd9, 5'd7, 1'd1} : fbdiv_cal_expected = 10'b0000011100;
  {SERDES, 4'd12, 5'd0, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd12, 5'd1, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd12, 5'd2, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd12, 5'd3, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd12, 5'd4, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd12, 5'd5, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd12, 5'd6, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd12, 5'd7, 1'd1} : fbdiv_cal_expected = 10'b0000010100;
  {SERDES, 4'd13, 5'd0, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd13, 5'd1, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd13, 5'd2, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd13, 5'd3, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd13, 5'd4, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd13, 5'd5, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd13, 5'd6, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SERDES, 4'd13, 5'd7, 1'd1} : fbdiv_cal_expected = 10'b0000010101;
  {SAS, 4'd0, 5'd0, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd0, 5'd1, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd0, 5'd2, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd0, 5'd3, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd0, 5'd4, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd0, 5'd5, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd0, 5'd6, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd0, 5'd7, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd1, 5'd0, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd1, 5'd1, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd1, 5'd2, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd1, 5'd3, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd1, 5'd4, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd1, 5'd5, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd1, 5'd6, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd1, 5'd7, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd2, 5'd0, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd2, 5'd1, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd2, 5'd2, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd2, 5'd3, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd2, 5'd4, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd2, 5'd5, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd2, 5'd6, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd2, 5'd7, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd3, 5'd0, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd3, 5'd1, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd3, 5'd2, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd3, 5'd3, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd3, 5'd4, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd3, 5'd5, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd3, 5'd6, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd3, 5'd7, 1'd1} : fbdiv_cal_expected = 10'b0000011000;
  {SAS, 4'd4, 5'd0, 1'd1} : fbdiv_cal_expected = 10'b0000010111;
  {SAS, 4'd4, 5'd1, 1'd1} : fbdiv_cal_expected = 10'b0000010111;
  {SAS, 4'd4, 5'd2, 1'd1} : fbdiv_cal_expected = 10'b0000010111;
  {SAS, 4'd4, 5'd3, 1'd1} : fbdiv_cal_expected = 10'b0000010111;
  {SAS, 4'd4, 5'd4, 1'd1} : fbdiv_cal_expected = 10'b0000010111;
  {SAS, 4'd4, 5'd5, 1'd1} : fbdiv_cal_expected = 10'b0000010111;
  {SAS, 4'd4, 5'd6, 1'd1} : fbdiv_cal_expected = 10'b0000010111;
  {SAS, 4'd4, 5'd7, 1'd1} : fbdiv_cal_expected = 10'b0000010111;
  {PCIE, 4'd2, 5'd0, 1'd1} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd2, 5'd1, 1'd1} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd2, 5'd2, 1'd1} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd2, 5'd3, 1'd1} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd2, 5'd4, 1'd1} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd2, 5'd5, 1'd1} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd2, 5'd6, 1'd1} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd2, 5'd7, 1'd1} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd3, 5'd0, 1'd1} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd3, 5'd1, 1'd1} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd3, 5'd2, 1'd1} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd3, 5'd3, 1'd1} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd3, 5'd4, 1'd1} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd3, 5'd5, 1'd1} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd3, 5'd6, 1'd1} : fbdiv_cal_expected = 10'b0000010000;
  {PCIE, 4'd3, 5'd7, 1'd1} : fbdiv_cal_expected = 10'b0000010000;
default: fbdiv_cal_expected = 10'bzzzzzzzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel} )
  {USB, 4'd1, 5'd0, 1'd0} : refdiv_expected = 4'b0001;
  {USB, 4'd1, 5'd1, 1'd0} : refdiv_expected = 4'b0001;
  {USB, 4'd1, 5'd2, 1'd0} : refdiv_expected = 4'b0001;
  {USB, 4'd1, 5'd3, 1'd0} : refdiv_expected = 4'b0001;
  {USB, 4'd1, 5'd4, 1'd0} : refdiv_expected = 4'b0001;
  {USB, 4'd1, 5'd5, 1'd0} : refdiv_expected = 4'b0010;
  {USB, 4'd1, 5'd6, 1'd0} : refdiv_expected = 4'b0001;
  {USB, 4'd1, 5'd7, 1'd0} : refdiv_expected = 4'b0010;
  {USB, 4'd2, 5'd0, 1'd0} : refdiv_expected = 4'b0001;
  {USB, 4'd2, 5'd1, 1'd0} : refdiv_expected = 4'b0001;
  {USB, 4'd2, 5'd2, 1'd0} : refdiv_expected = 4'b0001;
  {USB, 4'd2, 5'd3, 1'd0} : refdiv_expected = 4'b0001;
  {USB, 4'd2, 5'd4, 1'd0} : refdiv_expected = 4'b0001;
  {USB, 4'd2, 5'd5, 1'd0} : refdiv_expected = 4'b0010;
  {USB, 4'd2, 5'd6, 1'd0} : refdiv_expected = 4'b0001;
  {USB, 4'd2, 5'd7, 1'd0} : refdiv_expected = 4'b0010;
  {SERDES, 4'd0, 5'd0, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd0, 5'd1, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd0, 5'd2, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd0, 5'd3, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd0, 5'd4, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd0, 5'd5, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd0, 5'd6, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd0, 5'd7, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd1, 5'd0, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd1, 5'd1, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd1, 5'd2, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd1, 5'd3, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd1, 5'd4, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd1, 5'd5, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd1, 5'd6, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd1, 5'd7, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd2, 5'd0, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd2, 5'd1, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd2, 5'd2, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd2, 5'd3, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd2, 5'd4, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd2, 5'd5, 1'd0} : refdiv_expected = 4'b0010;
  {SERDES, 4'd2, 5'd6, 1'd0} : refdiv_expected = 4'b0010;
  {SERDES, 4'd2, 5'd7, 1'd0} : refdiv_expected = 4'b0010;
  {SERDES, 4'd3, 5'd0, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd3, 5'd1, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd3, 5'd2, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd3, 5'd3, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd3, 5'd4, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd3, 5'd5, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd3, 5'd6, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd3, 5'd7, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd4, 5'd0, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd4, 5'd1, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd4, 5'd2, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd4, 5'd3, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd4, 5'd4, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd4, 5'd5, 1'd0} : refdiv_expected = 4'b0010;
  {SERDES, 4'd4, 5'd6, 1'd0} : refdiv_expected = 4'b0010;
  {SERDES, 4'd4, 5'd7, 1'd0} : refdiv_expected = 4'b0010;
  {SERDES, 4'd5, 5'd0, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd5, 5'd1, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd5, 5'd2, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd5, 5'd3, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd5, 5'd4, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd5, 5'd5, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd5, 5'd6, 1'd0} : refdiv_expected = 4'b0010;
  {SERDES, 4'd5, 5'd7, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd6, 5'd0, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd6, 5'd1, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd6, 5'd2, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd6, 5'd3, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd6, 5'd4, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd6, 5'd5, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd6, 5'd6, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd6, 5'd7, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd7, 5'd0, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd7, 5'd1, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd7, 5'd2, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd7, 5'd3, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd7, 5'd4, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd7, 5'd5, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd7, 5'd6, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd7, 5'd7, 1'd0} : refdiv_expected = 4'b0010;
  {SERDES, 4'd8, 5'd0, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd8, 5'd1, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd8, 5'd2, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd8, 5'd3, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd8, 5'd4, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd8, 5'd5, 1'd0} : refdiv_expected = 4'b0010;
  {SERDES, 4'd8, 5'd6, 1'd0} : refdiv_expected = 4'b0010;
  {SERDES, 4'd8, 5'd7, 1'd0} : refdiv_expected = 4'b0010;
  {SERDES, 4'd9, 5'd0, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd9, 5'd1, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd9, 5'd2, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd9, 5'd3, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd9, 5'd4, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd9, 5'd5, 1'd0} : refdiv_expected = 4'b0010;
  {SERDES, 4'd9, 5'd6, 1'd0} : refdiv_expected = 4'b0010;
  {SERDES, 4'd9, 5'd7, 1'd0} : refdiv_expected = 4'b0010;
  {SERDES, 4'd12, 5'd0, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd12, 5'd1, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd12, 5'd2, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd12, 5'd3, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd12, 5'd4, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd12, 5'd5, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd12, 5'd6, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd12, 5'd7, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd13, 5'd0, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd13, 5'd1, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd13, 5'd2, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd13, 5'd3, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd13, 5'd4, 1'd0} : refdiv_expected = 4'b0001;
  {SERDES, 4'd13, 5'd5, 1'd0} : refdiv_expected = 4'b0010;
  {SERDES, 4'd13, 5'd6, 1'd0} : refdiv_expected = 4'b0010;
  {SERDES, 4'd13, 5'd7, 1'd0} : refdiv_expected = 4'b0010;
  {SAS, 4'd0, 5'd0, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd0, 5'd1, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd0, 5'd2, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd0, 5'd3, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd0, 5'd4, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd0, 5'd5, 1'd0} : refdiv_expected = 4'b0010;
  {SAS, 4'd0, 5'd6, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd0, 5'd7, 1'd0} : refdiv_expected = 4'b0100;
  {SAS, 4'd1, 5'd0, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd1, 5'd1, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd1, 5'd2, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd1, 5'd3, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd1, 5'd4, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd1, 5'd5, 1'd0} : refdiv_expected = 4'b0010;
  {SAS, 4'd1, 5'd6, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd1, 5'd7, 1'd0} : refdiv_expected = 4'b0100;
  {SAS, 4'd2, 5'd0, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd2, 5'd1, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd2, 5'd2, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd2, 5'd3, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd2, 5'd4, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd2, 5'd5, 1'd0} : refdiv_expected = 4'b0010;
  {SAS, 4'd2, 5'd6, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd2, 5'd7, 1'd0} : refdiv_expected = 4'b0100;
  {SAS, 4'd3, 5'd0, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd3, 5'd1, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd3, 5'd2, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd3, 5'd3, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd3, 5'd4, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd3, 5'd5, 1'd0} : refdiv_expected = 4'b0010;
  {SAS, 4'd3, 5'd6, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd3, 5'd7, 1'd0} : refdiv_expected = 4'b0100;
  {SAS, 4'd4, 5'd0, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd4, 5'd1, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd4, 5'd2, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd4, 5'd3, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd4, 5'd4, 1'd0} : refdiv_expected = 4'b0010;
  {SAS, 4'd4, 5'd5, 1'd0} : refdiv_expected = 4'b0010;
  {SAS, 4'd4, 5'd6, 1'd0} : refdiv_expected = 4'b0001;
  {SAS, 4'd4, 5'd7, 1'd0} : refdiv_expected = 4'b0010;
  {PCIE, 4'd2, 5'd0, 1'd0} : refdiv_expected = 4'b0001;
  {PCIE, 4'd2, 5'd1, 1'd0} : refdiv_expected = 4'b0001;
  {PCIE, 4'd2, 5'd2, 1'd0} : refdiv_expected = 4'b0001;
  {PCIE, 4'd2, 5'd3, 1'd0} : refdiv_expected = 4'b0010;
  {PCIE, 4'd2, 5'd4, 1'd0} : refdiv_expected = 4'b0001;
  {PCIE, 4'd2, 5'd5, 1'd0} : refdiv_expected = 4'b0001;
  {PCIE, 4'd2, 5'd6, 1'd0} : refdiv_expected = 4'b0001;
  {PCIE, 4'd2, 5'd7, 1'd0} : refdiv_expected = 4'b0100;
  {PCIE, 4'd3, 5'd0, 1'd0} : refdiv_expected = 4'b0001;
  {PCIE, 4'd3, 5'd1, 1'd0} : refdiv_expected = 4'b0001;
  {PCIE, 4'd3, 5'd2, 1'd0} : refdiv_expected = 4'b0001;
  {PCIE, 4'd3, 5'd3, 1'd0} : refdiv_expected = 4'b0010;
  {PCIE, 4'd3, 5'd4, 1'd0} : refdiv_expected = 4'b0001;
  {PCIE, 4'd3, 5'd5, 1'd0} : refdiv_expected = 4'b0001;
  {PCIE, 4'd3, 5'd6, 1'd0} : refdiv_expected = 4'b0001;
  {PCIE, 4'd3, 5'd7, 1'd0} : refdiv_expected = 4'b0100;
  {USB, 4'd1, 5'd0, 1'd1} : refdiv_expected = 4'b0001;
  {USB, 4'd1, 5'd1, 1'd1} : refdiv_expected = 4'b0001;
  {USB, 4'd1, 5'd2, 1'd1} : refdiv_expected = 4'b0010;
  {USB, 4'd1, 5'd3, 1'd1} : refdiv_expected = 4'b0001;
  {USB, 4'd1, 5'd4, 1'd1} : refdiv_expected = 4'b0001;
  {USB, 4'd1, 5'd5, 1'd1} : refdiv_expected = 4'b0010;
  {USB, 4'd1, 5'd6, 1'd1} : refdiv_expected = 4'b0001;
  {USB, 4'd1, 5'd7, 1'd1} : refdiv_expected = 4'b0010;
  {USB, 4'd2, 5'd0, 1'd1} : refdiv_expected = 4'b0001;
  {USB, 4'd2, 5'd1, 1'd1} : refdiv_expected = 4'b0001;
  {USB, 4'd2, 5'd2, 1'd1} : refdiv_expected = 4'b0010;
  {USB, 4'd2, 5'd3, 1'd1} : refdiv_expected = 4'b0001;
  {USB, 4'd2, 5'd4, 1'd1} : refdiv_expected = 4'b0001;
  {USB, 4'd2, 5'd5, 1'd1} : refdiv_expected = 4'b0010;
  {USB, 4'd2, 5'd6, 1'd1} : refdiv_expected = 4'b0001;
  {USB, 4'd2, 5'd7, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd0, 5'd0, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd0, 5'd1, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd0, 5'd2, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd0, 5'd3, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd0, 5'd4, 1'd1} : refdiv_expected = 4'b0011;
  {SERDES, 4'd0, 5'd5, 1'd1} : refdiv_expected = 4'b0011;
  {SERDES, 4'd0, 5'd6, 1'd1} : refdiv_expected = 4'b0011;
  {SERDES, 4'd0, 5'd7, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd1, 5'd0, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd1, 5'd1, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd1, 5'd2, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd1, 5'd3, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd1, 5'd4, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd1, 5'd5, 1'd1} : refdiv_expected = 4'b0011;
  {SERDES, 4'd1, 5'd6, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd1, 5'd7, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd2, 5'd0, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd2, 5'd1, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd2, 5'd2, 1'd1} : refdiv_expected = 4'b0011;
  {SERDES, 4'd2, 5'd3, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd2, 5'd4, 1'd1} : refdiv_expected = 4'b0100;
  {SERDES, 4'd2, 5'd5, 1'd1} : refdiv_expected = 4'b0100;
  {SERDES, 4'd2, 5'd6, 1'd1} : refdiv_expected = 4'b0011;
  {SERDES, 4'd2, 5'd7, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd3, 5'd0, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd3, 5'd1, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd3, 5'd2, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd3, 5'd3, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd3, 5'd4, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd3, 5'd5, 1'd1} : refdiv_expected = 4'b0011;
  {SERDES, 4'd3, 5'd6, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd3, 5'd7, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd4, 5'd0, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd4, 5'd1, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd4, 5'd2, 1'd1} : refdiv_expected = 4'b0011;
  {SERDES, 4'd4, 5'd3, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd4, 5'd4, 1'd1} : refdiv_expected = 4'b0100;
  {SERDES, 4'd4, 5'd5, 1'd1} : refdiv_expected = 4'b0100;
  {SERDES, 4'd4, 5'd6, 1'd1} : refdiv_expected = 4'b0011;
  {SERDES, 4'd4, 5'd7, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd5, 5'd0, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd5, 5'd1, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd5, 5'd2, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd5, 5'd3, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd5, 5'd4, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd5, 5'd5, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd5, 5'd6, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd5, 5'd7, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd6, 5'd0, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd6, 5'd1, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd6, 5'd2, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd6, 5'd3, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd6, 5'd4, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd6, 5'd5, 1'd1} : refdiv_expected = 4'b0011;
  {SERDES, 4'd6, 5'd6, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd6, 5'd7, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd7, 5'd0, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd7, 5'd1, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd7, 5'd2, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd7, 5'd3, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd7, 5'd4, 1'd1} : refdiv_expected = 4'b0011;
  {SERDES, 4'd7, 5'd5, 1'd1} : refdiv_expected = 4'b0011;
  {SERDES, 4'd7, 5'd6, 1'd1} : refdiv_expected = 4'b0101;
  {SERDES, 4'd7, 5'd7, 1'd1} : refdiv_expected = 4'b0011;
  {SERDES, 4'd8, 5'd0, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd8, 5'd1, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd8, 5'd2, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd8, 5'd3, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd8, 5'd4, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd8, 5'd5, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd8, 5'd6, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd8, 5'd7, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd9, 5'd0, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd9, 5'd1, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd9, 5'd2, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd9, 5'd3, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd9, 5'd4, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd9, 5'd5, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd9, 5'd6, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd9, 5'd7, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd12, 5'd0, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd12, 5'd1, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd12, 5'd2, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd12, 5'd3, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd12, 5'd4, 1'd1} : refdiv_expected = 4'b0011;
  {SERDES, 4'd12, 5'd5, 1'd1} : refdiv_expected = 4'b0011;
  {SERDES, 4'd12, 5'd6, 1'd1} : refdiv_expected = 4'b0011;
  {SERDES, 4'd12, 5'd7, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd13, 5'd0, 1'd1} : refdiv_expected = 4'b0001;
  {SERDES, 4'd13, 5'd1, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd13, 5'd2, 1'd1} : refdiv_expected = 4'b0011;
  {SERDES, 4'd13, 5'd3, 1'd1} : refdiv_expected = 4'b0010;
  {SERDES, 4'd13, 5'd4, 1'd1} : refdiv_expected = 4'b0100;
  {SERDES, 4'd13, 5'd5, 1'd1} : refdiv_expected = 4'b0100;
  {SERDES, 4'd13, 5'd6, 1'd1} : refdiv_expected = 4'b0011;
  {SERDES, 4'd13, 5'd7, 1'd1} : refdiv_expected = 4'b0010;
  {SAS, 4'd0, 5'd0, 1'd1} : refdiv_expected = 4'b0001;
  {SAS, 4'd0, 5'd1, 1'd1} : refdiv_expected = 4'b0001;
  {SAS, 4'd0, 5'd2, 1'd1} : refdiv_expected = 4'b0011;
  {SAS, 4'd0, 5'd3, 1'd1} : refdiv_expected = 4'b0011;
  {SAS, 4'd0, 5'd4, 1'd1} : refdiv_expected = 4'b0001;
  {SAS, 4'd0, 5'd5, 1'd1} : refdiv_expected = 4'b0010;
  {SAS, 4'd0, 5'd6, 1'd1} : refdiv_expected = 4'b0001;
  {SAS, 4'd0, 5'd7, 1'd1} : refdiv_expected = 4'b0100;
  {SAS, 4'd1, 5'd0, 1'd1} : refdiv_expected = 4'b0001;
  {SAS, 4'd1, 5'd1, 1'd1} : refdiv_expected = 4'b0001;
  {SAS, 4'd1, 5'd2, 1'd1} : refdiv_expected = 4'b0011;
  {SAS, 4'd1, 5'd3, 1'd1} : refdiv_expected = 4'b0011;
  {SAS, 4'd1, 5'd4, 1'd1} : refdiv_expected = 4'b0001;
  {SAS, 4'd1, 5'd5, 1'd1} : refdiv_expected = 4'b0010;
  {SAS, 4'd1, 5'd6, 1'd1} : refdiv_expected = 4'b0001;
  {SAS, 4'd1, 5'd7, 1'd1} : refdiv_expected = 4'b0100;
  {SAS, 4'd2, 5'd0, 1'd1} : refdiv_expected = 4'b0001;
  {SAS, 4'd2, 5'd1, 1'd1} : refdiv_expected = 4'b0001;
  {SAS, 4'd2, 5'd2, 1'd1} : refdiv_expected = 4'b0011;
  {SAS, 4'd2, 5'd3, 1'd1} : refdiv_expected = 4'b0011;
  {SAS, 4'd2, 5'd4, 1'd1} : refdiv_expected = 4'b0001;
  {SAS, 4'd2, 5'd5, 1'd1} : refdiv_expected = 4'b0010;
  {SAS, 4'd2, 5'd6, 1'd1} : refdiv_expected = 4'b0001;
  {SAS, 4'd2, 5'd7, 1'd1} : refdiv_expected = 4'b0100;
  {SAS, 4'd3, 5'd0, 1'd1} : refdiv_expected = 4'b0001;
  {SAS, 4'd3, 5'd1, 1'd1} : refdiv_expected = 4'b0001;
  {SAS, 4'd3, 5'd2, 1'd1} : refdiv_expected = 4'b0011;
  {SAS, 4'd3, 5'd3, 1'd1} : refdiv_expected = 4'b0011;
  {SAS, 4'd3, 5'd4, 1'd1} : refdiv_expected = 4'b0001;
  {SAS, 4'd3, 5'd5, 1'd1} : refdiv_expected = 4'b0010;
  {SAS, 4'd3, 5'd6, 1'd1} : refdiv_expected = 4'b0001;
  {SAS, 4'd3, 5'd7, 1'd1} : refdiv_expected = 4'b0100;
  {SAS, 4'd4, 5'd0, 1'd1} : refdiv_expected = 4'b0001;
  {SAS, 4'd4, 5'd1, 1'd1} : refdiv_expected = 4'b0001;
  {SAS, 4'd4, 5'd2, 1'd1} : refdiv_expected = 4'b0001;
  {SAS, 4'd4, 5'd3, 1'd1} : refdiv_expected = 4'b0001;
  {SAS, 4'd4, 5'd4, 1'd1} : refdiv_expected = 4'b0010;
  {SAS, 4'd4, 5'd5, 1'd1} : refdiv_expected = 4'b0010;
  {SAS, 4'd4, 5'd6, 1'd1} : refdiv_expected = 4'b0010;
  {SAS, 4'd4, 5'd7, 1'd1} : refdiv_expected = 4'b0010;
  {PCIE, 4'd2, 5'd0, 1'd1} : refdiv_expected = 4'b0001;
  {PCIE, 4'd2, 5'd1, 1'd1} : refdiv_expected = 4'b0010;
  {PCIE, 4'd2, 5'd2, 1'd1} : refdiv_expected = 4'b0001;
  {PCIE, 4'd2, 5'd3, 1'd1} : refdiv_expected = 4'b0010;
  {PCIE, 4'd2, 5'd4, 1'd1} : refdiv_expected = 4'b0001;
  {PCIE, 4'd2, 5'd5, 1'd1} : refdiv_expected = 4'b0001;
  {PCIE, 4'd2, 5'd6, 1'd1} : refdiv_expected = 4'b0001;
  {PCIE, 4'd2, 5'd7, 1'd1} : refdiv_expected = 4'b0100;
  {PCIE, 4'd3, 5'd0, 1'd1} : refdiv_expected = 4'b0001;
  {PCIE, 4'd3, 5'd1, 1'd1} : refdiv_expected = 4'b0010;
  {PCIE, 4'd3, 5'd2, 1'd1} : refdiv_expected = 4'b0001;
  {PCIE, 4'd3, 5'd3, 1'd1} : refdiv_expected = 4'b0010;
  {PCIE, 4'd3, 5'd4, 1'd1} : refdiv_expected = 4'b0001;
  {PCIE, 4'd3, 5'd5, 1'd1} : refdiv_expected = 4'b0001;
  {PCIE, 4'd3, 5'd6, 1'd1} : refdiv_expected = 4'b0001;
  {PCIE, 4'd3, 5'd7, 1'd1} : refdiv_expected = 4'b0100;
default: refdiv_expected = 4'bzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel} )
  {USB, 4'd1, 5'd0, 1'd0} : vind_band_sel_expected = 1'b0;
  {USB, 4'd1, 5'd1, 1'd0} : vind_band_sel_expected = 1'b0;
  {USB, 4'd1, 5'd2, 1'd0} : vind_band_sel_expected = 1'b0;
  {USB, 4'd1, 5'd3, 1'd0} : vind_band_sel_expected = 1'b0;
  {USB, 4'd1, 5'd4, 1'd0} : vind_band_sel_expected = 1'b0;
  {USB, 4'd1, 5'd5, 1'd0} : vind_band_sel_expected = 1'b0;
  {USB, 4'd1, 5'd6, 1'd0} : vind_band_sel_expected = 1'b0;
  {USB, 4'd1, 5'd7, 1'd0} : vind_band_sel_expected = 1'b0;
  {USB, 4'd2, 5'd0, 1'd0} : vind_band_sel_expected = 1'b0;
  {USB, 4'd2, 5'd1, 1'd0} : vind_band_sel_expected = 1'b0;
  {USB, 4'd2, 5'd2, 1'd0} : vind_band_sel_expected = 1'b0;
  {USB, 4'd2, 5'd3, 1'd0} : vind_band_sel_expected = 1'b0;
  {USB, 4'd2, 5'd4, 1'd0} : vind_band_sel_expected = 1'b0;
  {USB, 4'd2, 5'd5, 1'd0} : vind_band_sel_expected = 1'b0;
  {USB, 4'd2, 5'd6, 1'd0} : vind_band_sel_expected = 1'b0;
  {USB, 4'd2, 5'd7, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd0, 5'd0, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd0, 5'd1, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd0, 5'd2, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd0, 5'd3, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd0, 5'd4, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd0, 5'd5, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd0, 5'd6, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd0, 5'd7, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd1, 5'd0, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd1, 5'd1, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd1, 5'd2, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd1, 5'd3, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd1, 5'd4, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd1, 5'd5, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd1, 5'd6, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd1, 5'd7, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd2, 5'd0, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd2, 5'd1, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd2, 5'd2, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd2, 5'd3, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd2, 5'd4, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd2, 5'd5, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd2, 5'd6, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd2, 5'd7, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd3, 5'd0, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd3, 5'd1, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd3, 5'd2, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd3, 5'd3, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd3, 5'd4, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd3, 5'd5, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd3, 5'd6, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd3, 5'd7, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd4, 5'd0, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd4, 5'd1, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd4, 5'd2, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd4, 5'd3, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd4, 5'd4, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd4, 5'd5, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd4, 5'd6, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd4, 5'd7, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd5, 5'd0, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd5, 5'd1, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd5, 5'd2, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd5, 5'd3, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd5, 5'd4, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd5, 5'd5, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd5, 5'd6, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd5, 5'd7, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd6, 5'd0, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd6, 5'd1, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd6, 5'd2, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd6, 5'd3, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd6, 5'd4, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd6, 5'd5, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd6, 5'd6, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd6, 5'd7, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd7, 5'd0, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd7, 5'd1, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd7, 5'd2, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd7, 5'd3, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd7, 5'd4, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd7, 5'd5, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd7, 5'd6, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd7, 5'd7, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd8, 5'd0, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd8, 5'd1, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd8, 5'd2, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd8, 5'd3, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd8, 5'd4, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd8, 5'd5, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd8, 5'd6, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd8, 5'd7, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd9, 5'd0, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd9, 5'd1, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd9, 5'd2, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd9, 5'd3, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd9, 5'd4, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd9, 5'd5, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd9, 5'd6, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd9, 5'd7, 1'd0} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd12, 5'd0, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd12, 5'd1, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd12, 5'd2, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd12, 5'd3, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd12, 5'd4, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd12, 5'd5, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd12, 5'd6, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd12, 5'd7, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd13, 5'd0, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd13, 5'd1, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd13, 5'd2, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd13, 5'd3, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd13, 5'd4, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd13, 5'd5, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd13, 5'd6, 1'd0} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd13, 5'd7, 1'd0} : vind_band_sel_expected = 1'b0;
  {SAS, 4'd0, 5'd0, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd0, 5'd1, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd0, 5'd2, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd0, 5'd3, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd0, 5'd4, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd0, 5'd5, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd0, 5'd6, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd0, 5'd7, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd1, 5'd0, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd1, 5'd1, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd1, 5'd2, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd1, 5'd3, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd1, 5'd4, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd1, 5'd5, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd1, 5'd6, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd1, 5'd7, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd2, 5'd0, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd2, 5'd1, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd2, 5'd2, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd2, 5'd3, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd2, 5'd4, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd2, 5'd5, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd2, 5'd6, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd2, 5'd7, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd3, 5'd0, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd3, 5'd1, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd3, 5'd2, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd3, 5'd3, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd3, 5'd4, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd3, 5'd5, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd3, 5'd6, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd3, 5'd7, 1'd0} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd4, 5'd0, 1'd0} : vind_band_sel_expected = 1'b0;
  {SAS, 4'd4, 5'd1, 1'd0} : vind_band_sel_expected = 1'b0;
  {SAS, 4'd4, 5'd2, 1'd0} : vind_band_sel_expected = 1'b0;
  {SAS, 4'd4, 5'd3, 1'd0} : vind_band_sel_expected = 1'b0;
  {SAS, 4'd4, 5'd4, 1'd0} : vind_band_sel_expected = 1'b0;
  {SAS, 4'd4, 5'd5, 1'd0} : vind_band_sel_expected = 1'b0;
  {SAS, 4'd4, 5'd6, 1'd0} : vind_band_sel_expected = 1'b0;
  {SAS, 4'd4, 5'd7, 1'd0} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd2, 5'd0, 1'd0} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd2, 5'd1, 1'd0} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd2, 5'd2, 1'd0} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd2, 5'd3, 1'd0} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd2, 5'd4, 1'd0} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd2, 5'd5, 1'd0} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd2, 5'd6, 1'd0} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd2, 5'd7, 1'd0} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd3, 5'd0, 1'd0} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd3, 5'd1, 1'd0} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd3, 5'd2, 1'd0} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd3, 5'd3, 1'd0} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd3, 5'd4, 1'd0} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd3, 5'd5, 1'd0} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd3, 5'd6, 1'd0} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd3, 5'd7, 1'd0} : vind_band_sel_expected = 1'b0;
  {USB, 4'd1, 5'd0, 1'd1} : vind_band_sel_expected = 1'b0;
  {USB, 4'd1, 5'd1, 1'd1} : vind_band_sel_expected = 1'b0;
  {USB, 4'd1, 5'd2, 1'd1} : vind_band_sel_expected = 1'b0;
  {USB, 4'd1, 5'd3, 1'd1} : vind_band_sel_expected = 1'b0;
  {USB, 4'd1, 5'd4, 1'd1} : vind_band_sel_expected = 1'b0;
  {USB, 4'd1, 5'd5, 1'd1} : vind_band_sel_expected = 1'b0;
  {USB, 4'd1, 5'd6, 1'd1} : vind_band_sel_expected = 1'b0;
  {USB, 4'd1, 5'd7, 1'd1} : vind_band_sel_expected = 1'b0;
  {USB, 4'd2, 5'd0, 1'd1} : vind_band_sel_expected = 1'b0;
  {USB, 4'd2, 5'd1, 1'd1} : vind_band_sel_expected = 1'b0;
  {USB, 4'd2, 5'd2, 1'd1} : vind_band_sel_expected = 1'b0;
  {USB, 4'd2, 5'd3, 1'd1} : vind_band_sel_expected = 1'b0;
  {USB, 4'd2, 5'd4, 1'd1} : vind_band_sel_expected = 1'b0;
  {USB, 4'd2, 5'd5, 1'd1} : vind_band_sel_expected = 1'b0;
  {USB, 4'd2, 5'd6, 1'd1} : vind_band_sel_expected = 1'b0;
  {USB, 4'd2, 5'd7, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd0, 5'd0, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd0, 5'd1, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd0, 5'd2, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd0, 5'd3, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd0, 5'd4, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd0, 5'd5, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd0, 5'd6, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd0, 5'd7, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd1, 5'd0, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd1, 5'd1, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd1, 5'd2, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd1, 5'd3, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd1, 5'd4, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd1, 5'd5, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd1, 5'd6, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd1, 5'd7, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd2, 5'd0, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd2, 5'd1, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd2, 5'd2, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd2, 5'd3, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd2, 5'd4, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd2, 5'd5, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd2, 5'd6, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd2, 5'd7, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd3, 5'd0, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd3, 5'd1, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd3, 5'd2, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd3, 5'd3, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd3, 5'd4, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd3, 5'd5, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd3, 5'd6, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd3, 5'd7, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd4, 5'd0, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd4, 5'd1, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd4, 5'd2, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd4, 5'd3, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd4, 5'd4, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd4, 5'd5, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd4, 5'd6, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd4, 5'd7, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd5, 5'd0, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd5, 5'd1, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd5, 5'd2, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd5, 5'd3, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd5, 5'd4, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd5, 5'd5, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd5, 5'd6, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd5, 5'd7, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd6, 5'd0, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd6, 5'd1, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd6, 5'd2, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd6, 5'd3, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd6, 5'd4, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd6, 5'd5, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd6, 5'd6, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd6, 5'd7, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd7, 5'd0, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd7, 5'd1, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd7, 5'd2, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd7, 5'd3, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd7, 5'd4, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd7, 5'd5, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd7, 5'd6, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd7, 5'd7, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd8, 5'd0, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd8, 5'd1, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd8, 5'd2, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd8, 5'd3, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd8, 5'd4, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd8, 5'd5, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd8, 5'd6, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd8, 5'd7, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd9, 5'd0, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd9, 5'd1, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd9, 5'd2, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd9, 5'd3, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd9, 5'd4, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd9, 5'd5, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd9, 5'd6, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd9, 5'd7, 1'd1} : vind_band_sel_expected = 1'b1;
  {SERDES, 4'd12, 5'd0, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd12, 5'd1, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd12, 5'd2, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd12, 5'd3, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd12, 5'd4, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd12, 5'd5, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd12, 5'd6, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd12, 5'd7, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd13, 5'd0, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd13, 5'd1, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd13, 5'd2, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd13, 5'd3, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd13, 5'd4, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd13, 5'd5, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd13, 5'd6, 1'd1} : vind_band_sel_expected = 1'b0;
  {SERDES, 4'd13, 5'd7, 1'd1} : vind_band_sel_expected = 1'b0;
  {SAS, 4'd0, 5'd0, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd0, 5'd1, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd0, 5'd2, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd0, 5'd3, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd0, 5'd4, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd0, 5'd5, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd0, 5'd6, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd0, 5'd7, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd1, 5'd0, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd1, 5'd1, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd1, 5'd2, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd1, 5'd3, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd1, 5'd4, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd1, 5'd5, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd1, 5'd6, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd1, 5'd7, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd2, 5'd0, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd2, 5'd1, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd2, 5'd2, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd2, 5'd3, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd2, 5'd4, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd2, 5'd5, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd2, 5'd6, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd2, 5'd7, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd3, 5'd0, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd3, 5'd1, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd3, 5'd2, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd3, 5'd3, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd3, 5'd4, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd3, 5'd5, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd3, 5'd6, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd3, 5'd7, 1'd1} : vind_band_sel_expected = 1'b1;
  {SAS, 4'd4, 5'd0, 1'd1} : vind_band_sel_expected = 1'b0;
  {SAS, 4'd4, 5'd1, 1'd1} : vind_band_sel_expected = 1'b0;
  {SAS, 4'd4, 5'd2, 1'd1} : vind_band_sel_expected = 1'b0;
  {SAS, 4'd4, 5'd3, 1'd1} : vind_band_sel_expected = 1'b0;
  {SAS, 4'd4, 5'd4, 1'd1} : vind_band_sel_expected = 1'b0;
  {SAS, 4'd4, 5'd5, 1'd1} : vind_band_sel_expected = 1'b0;
  {SAS, 4'd4, 5'd6, 1'd1} : vind_band_sel_expected = 1'b0;
  {SAS, 4'd4, 5'd7, 1'd1} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd2, 5'd0, 1'd1} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd2, 5'd1, 1'd1} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd2, 5'd2, 1'd1} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd2, 5'd3, 1'd1} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd2, 5'd4, 1'd1} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd2, 5'd5, 1'd1} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd2, 5'd6, 1'd1} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd2, 5'd7, 1'd1} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd3, 5'd0, 1'd1} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd3, 5'd1, 1'd1} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd3, 5'd2, 1'd1} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd3, 5'd3, 1'd1} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd3, 5'd4, 1'd1} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd3, 5'd5, 1'd1} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd3, 5'd6, 1'd1} : vind_band_sel_expected = 1'b0;
  {PCIE, 4'd3, 5'd7, 1'd1} : vind_band_sel_expected = 1'b0;
default: vind_band_sel_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel} )
  {USB, 4'd1, 5'd0, 1'd0} : div_1g_expected = 10'b0000101000;
  {USB, 4'd1, 5'd1, 1'd0} : div_1g_expected = 10'b0000101000;
  {USB, 4'd1, 5'd2, 1'd0} : div_1g_expected = 10'b0000101000;
  {USB, 4'd1, 5'd3, 1'd0} : div_1g_expected = 10'b0000101000;
  {USB, 4'd1, 5'd4, 1'd0} : div_1g_expected = 10'b0000101000;
  {USB, 4'd1, 5'd5, 1'd0} : div_1g_expected = 10'b0000101000;
  {USB, 4'd1, 5'd6, 1'd0} : div_1g_expected = 10'b0000101000;
  {USB, 4'd1, 5'd7, 1'd0} : div_1g_expected = 10'b0000101000;
  {USB, 4'd2, 5'd0, 1'd0} : div_1g_expected = 10'b0000101000;
  {USB, 4'd2, 5'd1, 1'd0} : div_1g_expected = 10'b0000101000;
  {USB, 4'd2, 5'd2, 1'd0} : div_1g_expected = 10'b0000101000;
  {USB, 4'd2, 5'd3, 1'd0} : div_1g_expected = 10'b0000101000;
  {USB, 4'd2, 5'd4, 1'd0} : div_1g_expected = 10'b0000101000;
  {USB, 4'd2, 5'd5, 1'd0} : div_1g_expected = 10'b0000101000;
  {USB, 4'd2, 5'd6, 1'd0} : div_1g_expected = 10'b0000101000;
  {USB, 4'd2, 5'd7, 1'd0} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd0, 5'd0, 1'd0} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd0, 5'd1, 1'd0} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd0, 5'd2, 1'd0} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd0, 5'd3, 1'd0} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd0, 5'd4, 1'd0} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd0, 5'd5, 1'd0} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd0, 5'd6, 1'd0} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd0, 5'd7, 1'd0} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd1, 5'd0, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd1, 5'd1, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd1, 5'd2, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd1, 5'd3, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd1, 5'd4, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd1, 5'd5, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd1, 5'd6, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd1, 5'd7, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd2, 5'd0, 1'd0} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd2, 5'd1, 1'd0} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd2, 5'd2, 1'd0} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd2, 5'd3, 1'd0} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd2, 5'd4, 1'd0} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd2, 5'd5, 1'd0} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd2, 5'd6, 1'd0} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd2, 5'd7, 1'd0} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd3, 5'd0, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd3, 5'd1, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd3, 5'd2, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd3, 5'd3, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd3, 5'd4, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd3, 5'd5, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd3, 5'd6, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd3, 5'd7, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd4, 5'd0, 1'd0} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd4, 5'd1, 1'd0} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd4, 5'd2, 1'd0} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd4, 5'd3, 1'd0} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd4, 5'd4, 1'd0} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd4, 5'd5, 1'd0} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd4, 5'd6, 1'd0} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd4, 5'd7, 1'd0} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd5, 5'd0, 1'd0} : div_1g_expected = 10'b0000110001;
  {SERDES, 4'd5, 5'd1, 1'd0} : div_1g_expected = 10'b0000110001;
  {SERDES, 4'd5, 5'd2, 1'd0} : div_1g_expected = 10'b0000110001;
  {SERDES, 4'd5, 5'd3, 1'd0} : div_1g_expected = 10'b0000110001;
  {SERDES, 4'd5, 5'd4, 1'd0} : div_1g_expected = 10'b0000110001;
  {SERDES, 4'd5, 5'd5, 1'd0} : div_1g_expected = 10'b0000110001;
  {SERDES, 4'd5, 5'd6, 1'd0} : div_1g_expected = 10'b0000110001;
  {SERDES, 4'd5, 5'd7, 1'd0} : div_1g_expected = 10'b0000110001;
  {SERDES, 4'd6, 5'd0, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd6, 5'd1, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd6, 5'd2, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd6, 5'd3, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd6, 5'd4, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd6, 5'd5, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd6, 5'd6, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd6, 5'd7, 1'd0} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd7, 5'd0, 1'd0} : div_1g_expected = 10'b0000110100;
  {SERDES, 4'd7, 5'd1, 1'd0} : div_1g_expected = 10'b0000110100;
  {SERDES, 4'd7, 5'd2, 1'd0} : div_1g_expected = 10'b0000110100;
  {SERDES, 4'd7, 5'd3, 1'd0} : div_1g_expected = 10'b0000110100;
  {SERDES, 4'd7, 5'd4, 1'd0} : div_1g_expected = 10'b0000110100;
  {SERDES, 4'd7, 5'd5, 1'd0} : div_1g_expected = 10'b0000110100;
  {SERDES, 4'd7, 5'd6, 1'd0} : div_1g_expected = 10'b0000110100;
  {SERDES, 4'd7, 5'd7, 1'd0} : div_1g_expected = 10'b0000110100;
  {SERDES, 4'd8, 5'd0, 1'd0} : div_1g_expected = 10'b0000110111;
  {SERDES, 4'd8, 5'd1, 1'd0} : div_1g_expected = 10'b0000110111;
  {SERDES, 4'd8, 5'd2, 1'd0} : div_1g_expected = 10'b0000110111;
  {SERDES, 4'd8, 5'd3, 1'd0} : div_1g_expected = 10'b0000110111;
  {SERDES, 4'd8, 5'd4, 1'd0} : div_1g_expected = 10'b0000110111;
  {SERDES, 4'd8, 5'd5, 1'd0} : div_1g_expected = 10'b0000110111;
  {SERDES, 4'd8, 5'd6, 1'd0} : div_1g_expected = 10'b0000110111;
  {SERDES, 4'd8, 5'd7, 1'd0} : div_1g_expected = 10'b0000110111;
  {SERDES, 4'd9, 5'd0, 1'd0} : div_1g_expected = 10'b0000111000;
  {SERDES, 4'd9, 5'd1, 1'd0} : div_1g_expected = 10'b0000111000;
  {SERDES, 4'd9, 5'd2, 1'd0} : div_1g_expected = 10'b0000111000;
  {SERDES, 4'd9, 5'd3, 1'd0} : div_1g_expected = 10'b0000111000;
  {SERDES, 4'd9, 5'd4, 1'd0} : div_1g_expected = 10'b0000111000;
  {SERDES, 4'd9, 5'd5, 1'd0} : div_1g_expected = 10'b0000111000;
  {SERDES, 4'd9, 5'd6, 1'd0} : div_1g_expected = 10'b0000111000;
  {SERDES, 4'd9, 5'd7, 1'd0} : div_1g_expected = 10'b0000111000;
  {SERDES, 4'd12, 5'd0, 1'd0} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd12, 5'd1, 1'd0} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd12, 5'd2, 1'd0} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd12, 5'd3, 1'd0} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd12, 5'd4, 1'd0} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd12, 5'd5, 1'd0} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd12, 5'd6, 1'd0} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd12, 5'd7, 1'd0} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd13, 5'd0, 1'd0} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd13, 5'd1, 1'd0} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd13, 5'd2, 1'd0} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd13, 5'd3, 1'd0} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd13, 5'd4, 1'd0} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd13, 5'd5, 1'd0} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd13, 5'd6, 1'd0} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd13, 5'd7, 1'd0} : div_1g_expected = 10'b0000101001;
  {SAS, 4'd0, 5'd0, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd0, 5'd1, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd0, 5'd2, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd0, 5'd3, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd0, 5'd4, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd0, 5'd5, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd0, 5'd6, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd0, 5'd7, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd1, 5'd0, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd1, 5'd1, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd1, 5'd2, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd1, 5'd3, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd1, 5'd4, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd1, 5'd5, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd1, 5'd6, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd1, 5'd7, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd2, 5'd0, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd2, 5'd1, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd2, 5'd2, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd2, 5'd3, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd2, 5'd4, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd2, 5'd5, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd2, 5'd6, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd2, 5'd7, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd3, 5'd0, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd3, 5'd1, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd3, 5'd2, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd3, 5'd3, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd3, 5'd4, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd3, 5'd5, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd3, 5'd6, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd3, 5'd7, 1'd0} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd4, 5'd0, 1'd0} : div_1g_expected = 10'b0000101101;
  {SAS, 4'd4, 5'd1, 1'd0} : div_1g_expected = 10'b0000101101;
  {SAS, 4'd4, 5'd2, 1'd0} : div_1g_expected = 10'b0000101101;
  {SAS, 4'd4, 5'd3, 1'd0} : div_1g_expected = 10'b0000101101;
  {SAS, 4'd4, 5'd4, 1'd0} : div_1g_expected = 10'b0000101101;
  {SAS, 4'd4, 5'd5, 1'd0} : div_1g_expected = 10'b0000101101;
  {SAS, 4'd4, 5'd6, 1'd0} : div_1g_expected = 10'b0000101101;
  {SAS, 4'd4, 5'd7, 1'd0} : div_1g_expected = 10'b0000101101;
  {PCIE, 4'd2, 5'd0, 1'd0} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd2, 5'd1, 1'd0} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd2, 5'd2, 1'd0} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd2, 5'd3, 1'd0} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd2, 5'd4, 1'd0} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd2, 5'd5, 1'd0} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd2, 5'd6, 1'd0} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd2, 5'd7, 1'd0} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd3, 5'd0, 1'd0} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd3, 5'd1, 1'd0} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd3, 5'd2, 1'd0} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd3, 5'd3, 1'd0} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd3, 5'd4, 1'd0} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd3, 5'd5, 1'd0} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd3, 5'd6, 1'd0} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd3, 5'd7, 1'd0} : div_1g_expected = 10'b0000100000;
  {USB, 4'd1, 5'd0, 1'd1} : div_1g_expected = 10'b0000101000;
  {USB, 4'd1, 5'd1, 1'd1} : div_1g_expected = 10'b0000101000;
  {USB, 4'd1, 5'd2, 1'd1} : div_1g_expected = 10'b0000101000;
  {USB, 4'd1, 5'd3, 1'd1} : div_1g_expected = 10'b0000101000;
  {USB, 4'd1, 5'd4, 1'd1} : div_1g_expected = 10'b0000101000;
  {USB, 4'd1, 5'd5, 1'd1} : div_1g_expected = 10'b0000101000;
  {USB, 4'd1, 5'd6, 1'd1} : div_1g_expected = 10'b0000101000;
  {USB, 4'd1, 5'd7, 1'd1} : div_1g_expected = 10'b0000101000;
  {USB, 4'd2, 5'd0, 1'd1} : div_1g_expected = 10'b0000101000;
  {USB, 4'd2, 5'd1, 1'd1} : div_1g_expected = 10'b0000101000;
  {USB, 4'd2, 5'd2, 1'd1} : div_1g_expected = 10'b0000101000;
  {USB, 4'd2, 5'd3, 1'd1} : div_1g_expected = 10'b0000101000;
  {USB, 4'd2, 5'd4, 1'd1} : div_1g_expected = 10'b0000101000;
  {USB, 4'd2, 5'd5, 1'd1} : div_1g_expected = 10'b0000101000;
  {USB, 4'd2, 5'd6, 1'd1} : div_1g_expected = 10'b0000101000;
  {USB, 4'd2, 5'd7, 1'd1} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd0, 5'd0, 1'd1} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd0, 5'd1, 1'd1} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd0, 5'd2, 1'd1} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd0, 5'd3, 1'd1} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd0, 5'd4, 1'd1} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd0, 5'd5, 1'd1} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd0, 5'd6, 1'd1} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd0, 5'd7, 1'd1} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd1, 5'd0, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd1, 5'd1, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd1, 5'd2, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd1, 5'd3, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd1, 5'd4, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd1, 5'd5, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd1, 5'd6, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd1, 5'd7, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd2, 5'd0, 1'd1} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd2, 5'd1, 1'd1} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd2, 5'd2, 1'd1} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd2, 5'd3, 1'd1} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd2, 5'd4, 1'd1} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd2, 5'd5, 1'd1} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd2, 5'd6, 1'd1} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd2, 5'd7, 1'd1} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd3, 5'd0, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd3, 5'd1, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd3, 5'd2, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd3, 5'd3, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd3, 5'd4, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd3, 5'd5, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd3, 5'd6, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd3, 5'd7, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd4, 5'd0, 1'd1} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd4, 5'd1, 1'd1} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd4, 5'd2, 1'd1} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd4, 5'd3, 1'd1} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd4, 5'd4, 1'd1} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd4, 5'd5, 1'd1} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd4, 5'd6, 1'd1} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd4, 5'd7, 1'd1} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd5, 5'd0, 1'd1} : div_1g_expected = 10'b0000110001;
  {SERDES, 4'd5, 5'd1, 1'd1} : div_1g_expected = 10'b0000110001;
  {SERDES, 4'd5, 5'd2, 1'd1} : div_1g_expected = 10'b0000110001;
  {SERDES, 4'd5, 5'd3, 1'd1} : div_1g_expected = 10'b0000110001;
  {SERDES, 4'd5, 5'd4, 1'd1} : div_1g_expected = 10'b0000110001;
  {SERDES, 4'd5, 5'd5, 1'd1} : div_1g_expected = 10'b0000110001;
  {SERDES, 4'd5, 5'd6, 1'd1} : div_1g_expected = 10'b0000110001;
  {SERDES, 4'd5, 5'd7, 1'd1} : div_1g_expected = 10'b0000110001;
  {SERDES, 4'd6, 5'd0, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd6, 5'd1, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd6, 5'd2, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd6, 5'd3, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd6, 5'd4, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd6, 5'd5, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd6, 5'd6, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd6, 5'd7, 1'd1} : div_1g_expected = 10'b0000110010;
  {SERDES, 4'd7, 5'd0, 1'd1} : div_1g_expected = 10'b0000110100;
  {SERDES, 4'd7, 5'd1, 1'd1} : div_1g_expected = 10'b0000110100;
  {SERDES, 4'd7, 5'd2, 1'd1} : div_1g_expected = 10'b0000110100;
  {SERDES, 4'd7, 5'd3, 1'd1} : div_1g_expected = 10'b0000110100;
  {SERDES, 4'd7, 5'd4, 1'd1} : div_1g_expected = 10'b0000110100;
  {SERDES, 4'd7, 5'd5, 1'd1} : div_1g_expected = 10'b0000110100;
  {SERDES, 4'd7, 5'd6, 1'd1} : div_1g_expected = 10'b0000110100;
  {SERDES, 4'd7, 5'd7, 1'd1} : div_1g_expected = 10'b0000110100;
  {SERDES, 4'd8, 5'd0, 1'd1} : div_1g_expected = 10'b0000110111;
  {SERDES, 4'd8, 5'd1, 1'd1} : div_1g_expected = 10'b0000110111;
  {SERDES, 4'd8, 5'd2, 1'd1} : div_1g_expected = 10'b0000110111;
  {SERDES, 4'd8, 5'd3, 1'd1} : div_1g_expected = 10'b0000110111;
  {SERDES, 4'd8, 5'd4, 1'd1} : div_1g_expected = 10'b0000110111;
  {SERDES, 4'd8, 5'd5, 1'd1} : div_1g_expected = 10'b0000110111;
  {SERDES, 4'd8, 5'd6, 1'd1} : div_1g_expected = 10'b0000110111;
  {SERDES, 4'd8, 5'd7, 1'd1} : div_1g_expected = 10'b0000110111;
  {SERDES, 4'd9, 5'd0, 1'd1} : div_1g_expected = 10'b0000111000;
  {SERDES, 4'd9, 5'd1, 1'd1} : div_1g_expected = 10'b0000111000;
  {SERDES, 4'd9, 5'd2, 1'd1} : div_1g_expected = 10'b0000111000;
  {SERDES, 4'd9, 5'd3, 1'd1} : div_1g_expected = 10'b0000111000;
  {SERDES, 4'd9, 5'd4, 1'd1} : div_1g_expected = 10'b0000111000;
  {SERDES, 4'd9, 5'd5, 1'd1} : div_1g_expected = 10'b0000111000;
  {SERDES, 4'd9, 5'd6, 1'd1} : div_1g_expected = 10'b0000111000;
  {SERDES, 4'd9, 5'd7, 1'd1} : div_1g_expected = 10'b0000111000;
  {SERDES, 4'd12, 5'd0, 1'd1} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd12, 5'd1, 1'd1} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd12, 5'd2, 1'd1} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd12, 5'd3, 1'd1} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd12, 5'd4, 1'd1} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd12, 5'd5, 1'd1} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd12, 5'd6, 1'd1} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd12, 5'd7, 1'd1} : div_1g_expected = 10'b0000101000;
  {SERDES, 4'd13, 5'd0, 1'd1} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd13, 5'd1, 1'd1} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd13, 5'd2, 1'd1} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd13, 5'd3, 1'd1} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd13, 5'd4, 1'd1} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd13, 5'd5, 1'd1} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd13, 5'd6, 1'd1} : div_1g_expected = 10'b0000101001;
  {SERDES, 4'd13, 5'd7, 1'd1} : div_1g_expected = 10'b0000101001;
  {SAS, 4'd0, 5'd0, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd0, 5'd1, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd0, 5'd2, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd0, 5'd3, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd0, 5'd4, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd0, 5'd5, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd0, 5'd6, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd0, 5'd7, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd1, 5'd0, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd1, 5'd1, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd1, 5'd2, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd1, 5'd3, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd1, 5'd4, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd1, 5'd5, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd1, 5'd6, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd1, 5'd7, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd2, 5'd0, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd2, 5'd1, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd2, 5'd2, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd2, 5'd3, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd2, 5'd4, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd2, 5'd5, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd2, 5'd6, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd2, 5'd7, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd3, 5'd0, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd3, 5'd1, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd3, 5'd2, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd3, 5'd3, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd3, 5'd4, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd3, 5'd5, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd3, 5'd6, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd3, 5'd7, 1'd1} : div_1g_expected = 10'b0000110000;
  {SAS, 4'd4, 5'd0, 1'd1} : div_1g_expected = 10'b0000101101;
  {SAS, 4'd4, 5'd1, 1'd1} : div_1g_expected = 10'b0000101101;
  {SAS, 4'd4, 5'd2, 1'd1} : div_1g_expected = 10'b0000101101;
  {SAS, 4'd4, 5'd3, 1'd1} : div_1g_expected = 10'b0000101101;
  {SAS, 4'd4, 5'd4, 1'd1} : div_1g_expected = 10'b0000101101;
  {SAS, 4'd4, 5'd5, 1'd1} : div_1g_expected = 10'b0000101101;
  {SAS, 4'd4, 5'd6, 1'd1} : div_1g_expected = 10'b0000101101;
  {SAS, 4'd4, 5'd7, 1'd1} : div_1g_expected = 10'b0000101101;
  {PCIE, 4'd2, 5'd0, 1'd1} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd2, 5'd1, 1'd1} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd2, 5'd2, 1'd1} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd2, 5'd3, 1'd1} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd2, 5'd4, 1'd1} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd2, 5'd5, 1'd1} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd2, 5'd6, 1'd1} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd2, 5'd7, 1'd1} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd3, 5'd0, 1'd1} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd3, 5'd1, 1'd1} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd3, 5'd2, 1'd1} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd3, 5'd3, 1'd1} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd3, 5'd4, 1'd1} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd3, 5'd5, 1'd1} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd3, 5'd6, 1'd1} : div_1g_expected = 10'b0000100000;
  {PCIE, 4'd3, 5'd7, 1'd1} : div_1g_expected = 10'b0000100000;
default: div_1g_expected = 10'bzzzzzzzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel} )
  {USB, 4'd1, 5'd0, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd1, 5'd1, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd1, 5'd2, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd1, 5'd3, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd1, 5'd4, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd1, 5'd5, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd1, 5'd6, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd1, 5'd7, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd2, 5'd0, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd2, 5'd1, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd2, 5'd2, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd2, 5'd3, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd2, 5'd4, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd2, 5'd5, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd2, 5'd6, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd2, 5'd7, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd0, 5'd0, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd0, 5'd1, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd0, 5'd2, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd0, 5'd3, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd0, 5'd4, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd0, 5'd5, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd0, 5'd6, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd0, 5'd7, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd1, 5'd0, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd1, 5'd1, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd1, 5'd2, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd1, 5'd3, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd1, 5'd4, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd1, 5'd5, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd1, 5'd6, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd1, 5'd7, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd2, 5'd0, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd2, 5'd1, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd2, 5'd2, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd2, 5'd3, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd2, 5'd4, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd2, 5'd5, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd2, 5'd6, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd2, 5'd7, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd3, 5'd0, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd3, 5'd1, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd3, 5'd2, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd3, 5'd3, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd3, 5'd4, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd3, 5'd5, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd3, 5'd6, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd3, 5'd7, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd4, 5'd0, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd4, 5'd1, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd4, 5'd2, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd4, 5'd3, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd4, 5'd4, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd4, 5'd5, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd4, 5'd6, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd4, 5'd7, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd5, 5'd0, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SERDES, 4'd5, 5'd1, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SERDES, 4'd5, 5'd2, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SERDES, 4'd5, 5'd3, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SERDES, 4'd5, 5'd4, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SERDES, 4'd5, 5'd5, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SERDES, 4'd5, 5'd6, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SERDES, 4'd5, 5'd7, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SERDES, 4'd6, 5'd0, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd6, 5'd1, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd6, 5'd2, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd6, 5'd3, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd6, 5'd4, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd6, 5'd5, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd6, 5'd6, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd6, 5'd7, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd7, 5'd0, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd7, 5'd1, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd7, 5'd2, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd7, 5'd3, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd7, 5'd4, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd7, 5'd5, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd7, 5'd6, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd7, 5'd7, 1'd0} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd8, 5'd0, 1'd0} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd8, 5'd1, 1'd0} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd8, 5'd2, 1'd0} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd8, 5'd3, 1'd0} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd8, 5'd4, 1'd0} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd8, 5'd5, 1'd0} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd8, 5'd6, 1'd0} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd8, 5'd7, 1'd0} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd9, 5'd0, 1'd0} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd9, 5'd1, 1'd0} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd9, 5'd2, 1'd0} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd9, 5'd3, 1'd0} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd9, 5'd4, 1'd0} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd9, 5'd5, 1'd0} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd9, 5'd6, 1'd0} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd9, 5'd7, 1'd0} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd12, 5'd0, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd12, 5'd1, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd12, 5'd2, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd12, 5'd3, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd12, 5'd4, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd12, 5'd5, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd12, 5'd6, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd12, 5'd7, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd13, 5'd0, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd13, 5'd1, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd13, 5'd2, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd13, 5'd3, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd13, 5'd4, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd13, 5'd5, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd13, 5'd6, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd13, 5'd7, 1'd0} : div_1g_fbck_expected = 10'b0000001010;
  {SAS, 4'd0, 5'd0, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd0, 5'd1, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd0, 5'd2, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd0, 5'd3, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd0, 5'd4, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd0, 5'd5, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd0, 5'd6, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd0, 5'd7, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd1, 5'd0, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd1, 5'd1, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd1, 5'd2, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd1, 5'd3, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd1, 5'd4, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd1, 5'd5, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd1, 5'd6, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd1, 5'd7, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd2, 5'd0, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd2, 5'd1, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd2, 5'd2, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd2, 5'd3, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd2, 5'd4, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd2, 5'd5, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd2, 5'd6, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd2, 5'd7, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd3, 5'd0, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd3, 5'd1, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd3, 5'd2, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd3, 5'd3, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd3, 5'd4, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd3, 5'd5, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd3, 5'd6, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd3, 5'd7, 1'd0} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd4, 5'd0, 1'd0} : div_1g_fbck_expected = 10'b0000001011;
  {SAS, 4'd4, 5'd1, 1'd0} : div_1g_fbck_expected = 10'b0000001011;
  {SAS, 4'd4, 5'd2, 1'd0} : div_1g_fbck_expected = 10'b0000001011;
  {SAS, 4'd4, 5'd3, 1'd0} : div_1g_fbck_expected = 10'b0000001011;
  {SAS, 4'd4, 5'd4, 1'd0} : div_1g_fbck_expected = 10'b0000001011;
  {SAS, 4'd4, 5'd5, 1'd0} : div_1g_fbck_expected = 10'b0000001011;
  {SAS, 4'd4, 5'd6, 1'd0} : div_1g_fbck_expected = 10'b0000001011;
  {SAS, 4'd4, 5'd7, 1'd0} : div_1g_fbck_expected = 10'b0000001011;
  {PCIE, 4'd2, 5'd0, 1'd0} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd2, 5'd1, 1'd0} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd2, 5'd2, 1'd0} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd2, 5'd3, 1'd0} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd2, 5'd4, 1'd0} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd2, 5'd5, 1'd0} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd2, 5'd6, 1'd0} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd2, 5'd7, 1'd0} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd3, 5'd0, 1'd0} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd3, 5'd1, 1'd0} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd3, 5'd2, 1'd0} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd3, 5'd3, 1'd0} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd3, 5'd4, 1'd0} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd3, 5'd5, 1'd0} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd3, 5'd6, 1'd0} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd3, 5'd7, 1'd0} : div_1g_fbck_expected = 10'b0000001000;
  {USB, 4'd1, 5'd0, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd1, 5'd1, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd1, 5'd2, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd1, 5'd3, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd1, 5'd4, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd1, 5'd5, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd1, 5'd6, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd1, 5'd7, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd2, 5'd0, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd2, 5'd1, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd2, 5'd2, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd2, 5'd3, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd2, 5'd4, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd2, 5'd5, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd2, 5'd6, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {USB, 4'd2, 5'd7, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd0, 5'd0, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd0, 5'd1, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd0, 5'd2, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd0, 5'd3, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd0, 5'd4, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd0, 5'd5, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd0, 5'd6, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd0, 5'd7, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd1, 5'd0, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd1, 5'd1, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd1, 5'd2, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd1, 5'd3, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd1, 5'd4, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd1, 5'd5, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd1, 5'd6, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd1, 5'd7, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd2, 5'd0, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd2, 5'd1, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd2, 5'd2, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd2, 5'd3, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd2, 5'd4, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd2, 5'd5, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd2, 5'd6, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd2, 5'd7, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd3, 5'd0, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd3, 5'd1, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd3, 5'd2, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd3, 5'd3, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd3, 5'd4, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd3, 5'd5, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd3, 5'd6, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd3, 5'd7, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd4, 5'd0, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd4, 5'd1, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd4, 5'd2, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd4, 5'd3, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd4, 5'd4, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd4, 5'd5, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd4, 5'd6, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd4, 5'd7, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd5, 5'd0, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SERDES, 4'd5, 5'd1, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SERDES, 4'd5, 5'd2, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SERDES, 4'd5, 5'd3, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SERDES, 4'd5, 5'd4, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SERDES, 4'd5, 5'd5, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SERDES, 4'd5, 5'd6, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SERDES, 4'd5, 5'd7, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SERDES, 4'd6, 5'd0, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd6, 5'd1, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd6, 5'd2, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd6, 5'd3, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd6, 5'd4, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd6, 5'd5, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd6, 5'd6, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd6, 5'd7, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd7, 5'd0, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd7, 5'd1, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd7, 5'd2, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd7, 5'd3, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd7, 5'd4, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd7, 5'd5, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd7, 5'd6, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd7, 5'd7, 1'd1} : div_1g_fbck_expected = 10'b0000001101;
  {SERDES, 4'd8, 5'd0, 1'd1} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd8, 5'd1, 1'd1} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd8, 5'd2, 1'd1} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd8, 5'd3, 1'd1} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd8, 5'd4, 1'd1} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd8, 5'd5, 1'd1} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd8, 5'd6, 1'd1} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd8, 5'd7, 1'd1} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd9, 5'd0, 1'd1} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd9, 5'd1, 1'd1} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd9, 5'd2, 1'd1} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd9, 5'd3, 1'd1} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd9, 5'd4, 1'd1} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd9, 5'd5, 1'd1} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd9, 5'd6, 1'd1} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd9, 5'd7, 1'd1} : div_1g_fbck_expected = 10'b0000001110;
  {SERDES, 4'd12, 5'd0, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd12, 5'd1, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd12, 5'd2, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd12, 5'd3, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd12, 5'd4, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd12, 5'd5, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd12, 5'd6, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd12, 5'd7, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd13, 5'd0, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd13, 5'd1, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd13, 5'd2, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd13, 5'd3, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd13, 5'd4, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd13, 5'd5, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd13, 5'd6, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SERDES, 4'd13, 5'd7, 1'd1} : div_1g_fbck_expected = 10'b0000001010;
  {SAS, 4'd0, 5'd0, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd0, 5'd1, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd0, 5'd2, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd0, 5'd3, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd0, 5'd4, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd0, 5'd5, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd0, 5'd6, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd0, 5'd7, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd1, 5'd0, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd1, 5'd1, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd1, 5'd2, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd1, 5'd3, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd1, 5'd4, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd1, 5'd5, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd1, 5'd6, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd1, 5'd7, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd2, 5'd0, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd2, 5'd1, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd2, 5'd2, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd2, 5'd3, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd2, 5'd4, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd2, 5'd5, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd2, 5'd6, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd2, 5'd7, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd3, 5'd0, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd3, 5'd1, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd3, 5'd2, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd3, 5'd3, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd3, 5'd4, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd3, 5'd5, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd3, 5'd6, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd3, 5'd7, 1'd1} : div_1g_fbck_expected = 10'b0000001100;
  {SAS, 4'd4, 5'd0, 1'd1} : div_1g_fbck_expected = 10'b0000001011;
  {SAS, 4'd4, 5'd1, 1'd1} : div_1g_fbck_expected = 10'b0000001011;
  {SAS, 4'd4, 5'd2, 1'd1} : div_1g_fbck_expected = 10'b0000001011;
  {SAS, 4'd4, 5'd3, 1'd1} : div_1g_fbck_expected = 10'b0000001011;
  {SAS, 4'd4, 5'd4, 1'd1} : div_1g_fbck_expected = 10'b0000001011;
  {SAS, 4'd4, 5'd5, 1'd1} : div_1g_fbck_expected = 10'b0000001011;
  {SAS, 4'd4, 5'd6, 1'd1} : div_1g_fbck_expected = 10'b0000001011;
  {SAS, 4'd4, 5'd7, 1'd1} : div_1g_fbck_expected = 10'b0000001011;
  {PCIE, 4'd2, 5'd0, 1'd1} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd2, 5'd1, 1'd1} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd2, 5'd2, 1'd1} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd2, 5'd3, 1'd1} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd2, 5'd4, 1'd1} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd2, 5'd5, 1'd1} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd2, 5'd6, 1'd1} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd2, 5'd7, 1'd1} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd3, 5'd0, 1'd1} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd3, 5'd1, 1'd1} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd3, 5'd2, 1'd1} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd3, 5'd3, 1'd1} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd3, 5'd4, 1'd1} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd3, 5'd5, 1'd1} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd3, 5'd6, 1'd1} : div_1g_fbck_expected = 10'b0000001000;
  {PCIE, 4'd3, 5'd7, 1'd1} : div_1g_fbck_expected = 10'b0000001000;
default: div_1g_fbck_expected = 10'bzzzzzzzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel} )
  {USB, 4'd1, 5'd0, 1'd0} : icp_lc_expected = 5'b01111;
  {USB, 4'd1, 5'd1, 1'd0} : icp_lc_expected = 5'b01111;
  {USB, 4'd1, 5'd2, 1'd0} : icp_lc_expected = 5'b01110;
  {USB, 4'd1, 5'd3, 1'd0} : icp_lc_expected = 5'b01101;
  {USB, 4'd1, 5'd4, 1'd0} : icp_lc_expected = 5'b01100;
  {USB, 4'd1, 5'd5, 1'd0} : icp_lc_expected = 5'b01101;
  {USB, 4'd1, 5'd6, 1'd0} : icp_lc_expected = 5'b01010;
  {USB, 4'd1, 5'd7, 1'd0} : icp_lc_expected = 5'b01100;
  {USB, 4'd2, 5'd0, 1'd0} : icp_lc_expected = 5'b01111;
  {USB, 4'd2, 5'd1, 1'd0} : icp_lc_expected = 5'b01111;
  {USB, 4'd2, 5'd2, 1'd0} : icp_lc_expected = 5'b01110;
  {USB, 4'd2, 5'd3, 1'd0} : icp_lc_expected = 5'b01101;
  {USB, 4'd2, 5'd4, 1'd0} : icp_lc_expected = 5'b01100;
  {USB, 4'd2, 5'd5, 1'd0} : icp_lc_expected = 5'b01101;
  {USB, 4'd2, 5'd6, 1'd0} : icp_lc_expected = 5'b01010;
  {USB, 4'd2, 5'd7, 1'd0} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd0, 5'd0, 1'd0} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd0, 5'd1, 1'd0} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd0, 5'd2, 1'd0} : icp_lc_expected = 5'b01101;
  {SERDES, 4'd0, 5'd3, 1'd0} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd0, 5'd4, 1'd0} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd0, 5'd5, 1'd0} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd0, 5'd6, 1'd0} : icp_lc_expected = 5'b01010;
  {SERDES, 4'd0, 5'd7, 1'd0} : icp_lc_expected = 5'b01001;
  {SERDES, 4'd1, 5'd0, 1'd0} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd1, 5'd1, 1'd0} : icp_lc_expected = 5'b01101;
  {SERDES, 4'd1, 5'd2, 1'd0} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd1, 5'd3, 1'd0} : icp_lc_expected = 5'b01010;
  {SERDES, 4'd1, 5'd4, 1'd0} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd1, 5'd5, 1'd0} : icp_lc_expected = 5'b01000;
  {SERDES, 4'd1, 5'd6, 1'd0} : icp_lc_expected = 5'b00111;
  {SERDES, 4'd1, 5'd7, 1'd0} : icp_lc_expected = 5'b00110;
  {SERDES, 4'd2, 5'd0, 1'd0} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd2, 5'd1, 1'd0} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd2, 5'd2, 1'd0} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd2, 5'd3, 1'd0} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd2, 5'd4, 1'd0} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd2, 5'd5, 1'd0} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd2, 5'd6, 1'd0} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd2, 5'd7, 1'd0} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd3, 5'd0, 1'd0} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd3, 5'd1, 1'd0} : icp_lc_expected = 5'b01101;
  {SERDES, 4'd3, 5'd2, 1'd0} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd3, 5'd3, 1'd0} : icp_lc_expected = 5'b01010;
  {SERDES, 4'd3, 5'd4, 1'd0} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd3, 5'd5, 1'd0} : icp_lc_expected = 5'b01000;
  {SERDES, 4'd3, 5'd6, 1'd0} : icp_lc_expected = 5'b00111;
  {SERDES, 4'd3, 5'd7, 1'd0} : icp_lc_expected = 5'b00110;
  {SERDES, 4'd4, 5'd0, 1'd0} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd4, 5'd1, 1'd0} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd4, 5'd2, 1'd0} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd4, 5'd3, 1'd0} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd4, 5'd4, 1'd0} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd4, 5'd5, 1'd0} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd4, 5'd6, 1'd0} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd4, 5'd7, 1'd0} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd5, 5'd0, 1'd0} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd5, 5'd1, 1'd0} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd5, 5'd2, 1'd0} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd5, 5'd3, 1'd0} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd5, 5'd4, 1'd0} : icp_lc_expected = 5'b01101;
  {SERDES, 4'd5, 5'd5, 1'd0} : icp_lc_expected = 5'b01010;
  {SERDES, 4'd5, 5'd6, 1'd0} : icp_lc_expected = 5'b01101;
  {SERDES, 4'd5, 5'd7, 1'd0} : icp_lc_expected = 5'b01000;
  {SERDES, 4'd6, 5'd0, 1'd0} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd6, 5'd1, 1'd0} : icp_lc_expected = 5'b01101;
  {SERDES, 4'd6, 5'd2, 1'd0} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd6, 5'd3, 1'd0} : icp_lc_expected = 5'b01010;
  {SERDES, 4'd6, 5'd4, 1'd0} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd6, 5'd5, 1'd0} : icp_lc_expected = 5'b01000;
  {SERDES, 4'd6, 5'd6, 1'd0} : icp_lc_expected = 5'b00111;
  {SERDES, 4'd6, 5'd7, 1'd0} : icp_lc_expected = 5'b00110;
  {SERDES, 4'd7, 5'd0, 1'd0} : icp_lc_expected = 5'b01101;
  {SERDES, 4'd7, 5'd1, 1'd0} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd7, 5'd2, 1'd0} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd7, 5'd3, 1'd0} : icp_lc_expected = 5'b01010;
  {SERDES, 4'd7, 5'd4, 1'd0} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd7, 5'd5, 1'd0} : icp_lc_expected = 5'b01000;
  {SERDES, 4'd7, 5'd6, 1'd0} : icp_lc_expected = 5'b00111;
  {SERDES, 4'd7, 5'd7, 1'd0} : icp_lc_expected = 5'b01001;
  {SERDES, 4'd8, 5'd0, 1'd0} : icp_lc_expected = 5'b01101;
  {SERDES, 4'd8, 5'd1, 1'd0} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd8, 5'd2, 1'd0} : icp_lc_expected = 5'b01010;
  {SERDES, 4'd8, 5'd3, 1'd0} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd8, 5'd4, 1'd0} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd8, 5'd5, 1'd0} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd8, 5'd6, 1'd0} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd8, 5'd7, 1'd0} : icp_lc_expected = 5'b01001;
  {SERDES, 4'd9, 5'd0, 1'd0} : icp_lc_expected = 5'b01101;
  {SERDES, 4'd9, 5'd1, 1'd0} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd9, 5'd2, 1'd0} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd9, 5'd3, 1'd0} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd9, 5'd4, 1'd0} : icp_lc_expected = 5'b01010;
  {SERDES, 4'd9, 5'd5, 1'd0} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd9, 5'd6, 1'd0} : icp_lc_expected = 5'b01010;
  {SERDES, 4'd9, 5'd7, 1'd0} : icp_lc_expected = 5'b01001;
  {SERDES, 4'd12, 5'd0, 1'd0} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd12, 5'd1, 1'd0} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd12, 5'd2, 1'd0} : icp_lc_expected = 5'b01101;
  {SERDES, 4'd12, 5'd3, 1'd0} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd12, 5'd4, 1'd0} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd12, 5'd5, 1'd0} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd12, 5'd6, 1'd0} : icp_lc_expected = 5'b01010;
  {SERDES, 4'd12, 5'd7, 1'd0} : icp_lc_expected = 5'b01001;
  {SERDES, 4'd13, 5'd0, 1'd0} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd13, 5'd1, 1'd0} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd13, 5'd2, 1'd0} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd13, 5'd3, 1'd0} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd13, 5'd4, 1'd0} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd13, 5'd5, 1'd0} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd13, 5'd6, 1'd0} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd13, 5'd7, 1'd0} : icp_lc_expected = 5'b01100;
  {SAS, 4'd0, 5'd0, 1'd0} : icp_lc_expected = 5'b01111;
  {SAS, 4'd0, 5'd1, 1'd0} : icp_lc_expected = 5'b01111;
  {SAS, 4'd0, 5'd2, 1'd0} : icp_lc_expected = 5'b01101;
  {SAS, 4'd0, 5'd3, 1'd0} : icp_lc_expected = 5'b01100;
  {SAS, 4'd0, 5'd4, 1'd0} : icp_lc_expected = 5'b01010;
  {SAS, 4'd0, 5'd5, 1'd0} : icp_lc_expected = 5'b01100;
  {SAS, 4'd0, 5'd6, 1'd0} : icp_lc_expected = 5'b01001;
  {SAS, 4'd0, 5'd7, 1'd0} : icp_lc_expected = 5'b01101;
  {SAS, 4'd1, 5'd0, 1'd0} : icp_lc_expected = 5'b01111;
  {SAS, 4'd1, 5'd1, 1'd0} : icp_lc_expected = 5'b01111;
  {SAS, 4'd1, 5'd2, 1'd0} : icp_lc_expected = 5'b01101;
  {SAS, 4'd1, 5'd3, 1'd0} : icp_lc_expected = 5'b01100;
  {SAS, 4'd1, 5'd4, 1'd0} : icp_lc_expected = 5'b01010;
  {SAS, 4'd1, 5'd5, 1'd0} : icp_lc_expected = 5'b01100;
  {SAS, 4'd1, 5'd6, 1'd0} : icp_lc_expected = 5'b01001;
  {SAS, 4'd1, 5'd7, 1'd0} : icp_lc_expected = 5'b01101;
  {SAS, 4'd2, 5'd0, 1'd0} : icp_lc_expected = 5'b01111;
  {SAS, 4'd2, 5'd1, 1'd0} : icp_lc_expected = 5'b01111;
  {SAS, 4'd2, 5'd2, 1'd0} : icp_lc_expected = 5'b01101;
  {SAS, 4'd2, 5'd3, 1'd0} : icp_lc_expected = 5'b01100;
  {SAS, 4'd2, 5'd4, 1'd0} : icp_lc_expected = 5'b01010;
  {SAS, 4'd2, 5'd5, 1'd0} : icp_lc_expected = 5'b01100;
  {SAS, 4'd2, 5'd6, 1'd0} : icp_lc_expected = 5'b01001;
  {SAS, 4'd2, 5'd7, 1'd0} : icp_lc_expected = 5'b01101;
  {SAS, 4'd3, 5'd0, 1'd0} : icp_lc_expected = 5'b01111;
  {SAS, 4'd3, 5'd1, 1'd0} : icp_lc_expected = 5'b01111;
  {SAS, 4'd3, 5'd2, 1'd0} : icp_lc_expected = 5'b01101;
  {SAS, 4'd3, 5'd3, 1'd0} : icp_lc_expected = 5'b01100;
  {SAS, 4'd3, 5'd4, 1'd0} : icp_lc_expected = 5'b01010;
  {SAS, 4'd3, 5'd5, 1'd0} : icp_lc_expected = 5'b01100;
  {SAS, 4'd3, 5'd6, 1'd0} : icp_lc_expected = 5'b01001;
  {SAS, 4'd3, 5'd7, 1'd0} : icp_lc_expected = 5'b01101;
  {SAS, 4'd4, 5'd0, 1'd0} : icp_lc_expected = 5'b01111;
  {SAS, 4'd4, 5'd1, 1'd0} : icp_lc_expected = 5'b01111;
  {SAS, 4'd4, 5'd2, 1'd0} : icp_lc_expected = 5'b01101;
  {SAS, 4'd4, 5'd3, 1'd0} : icp_lc_expected = 5'b01100;
  {SAS, 4'd4, 5'd4, 1'd0} : icp_lc_expected = 5'b01110;
  {SAS, 4'd4, 5'd5, 1'd0} : icp_lc_expected = 5'b01100;
  {SAS, 4'd4, 5'd6, 1'd0} : icp_lc_expected = 5'b01001;
  {SAS, 4'd4, 5'd7, 1'd0} : icp_lc_expected = 5'b01100;
  {PCIE, 4'd2, 5'd0, 1'd0} : icp_lc_expected = 5'b01111;
  {PCIE, 4'd2, 5'd1, 1'd0} : icp_lc_expected = 5'b01111;
  {PCIE, 4'd2, 5'd2, 1'd0} : icp_lc_expected = 5'b01111;
  {PCIE, 4'd2, 5'd3, 1'd0} : icp_lc_expected = 5'b01111;
  {PCIE, 4'd2, 5'd4, 1'd0} : icp_lc_expected = 5'b01101;
  {PCIE, 4'd2, 5'd5, 1'd0} : icp_lc_expected = 5'b01111;
  {PCIE, 4'd2, 5'd6, 1'd0} : icp_lc_expected = 5'b01011;
  {PCIE, 4'd2, 5'd7, 1'd0} : icp_lc_expected = 5'b01111;
  {PCIE, 4'd3, 5'd0, 1'd0} : icp_lc_expected = 5'b01111;
  {PCIE, 4'd3, 5'd1, 1'd0} : icp_lc_expected = 5'b01111;
  {PCIE, 4'd3, 5'd2, 1'd0} : icp_lc_expected = 5'b01111;
  {PCIE, 4'd3, 5'd3, 1'd0} : icp_lc_expected = 5'b01111;
  {PCIE, 4'd3, 5'd4, 1'd0} : icp_lc_expected = 5'b01101;
  {PCIE, 4'd3, 5'd5, 1'd0} : icp_lc_expected = 5'b01111;
  {PCIE, 4'd3, 5'd6, 1'd0} : icp_lc_expected = 5'b01011;
  {PCIE, 4'd3, 5'd7, 1'd0} : icp_lc_expected = 5'b01111;
  {USB, 4'd1, 5'd0, 1'd1} : icp_lc_expected = 5'b01111;
  {USB, 4'd1, 5'd1, 1'd1} : icp_lc_expected = 5'b01111;
  {USB, 4'd1, 5'd2, 1'd1} : icp_lc_expected = 5'b01111;
  {USB, 4'd1, 5'd3, 1'd1} : icp_lc_expected = 5'b01101;
  {USB, 4'd1, 5'd4, 1'd1} : icp_lc_expected = 5'b01100;
  {USB, 4'd1, 5'd5, 1'd1} : icp_lc_expected = 5'b01101;
  {USB, 4'd1, 5'd6, 1'd1} : icp_lc_expected = 5'b01010;
  {USB, 4'd1, 5'd7, 1'd1} : icp_lc_expected = 5'b01100;
  {USB, 4'd2, 5'd0, 1'd1} : icp_lc_expected = 5'b01111;
  {USB, 4'd2, 5'd1, 1'd1} : icp_lc_expected = 5'b01111;
  {USB, 4'd2, 5'd2, 1'd1} : icp_lc_expected = 5'b01111;
  {USB, 4'd2, 5'd3, 1'd1} : icp_lc_expected = 5'b01101;
  {USB, 4'd2, 5'd4, 1'd1} : icp_lc_expected = 5'b01100;
  {USB, 4'd2, 5'd5, 1'd1} : icp_lc_expected = 5'b01101;
  {USB, 4'd2, 5'd6, 1'd1} : icp_lc_expected = 5'b01010;
  {USB, 4'd2, 5'd7, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd0, 5'd0, 1'd1} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd0, 5'd1, 1'd1} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd0, 5'd2, 1'd1} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd0, 5'd3, 1'd1} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd0, 5'd4, 1'd1} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd0, 5'd5, 1'd1} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd0, 5'd6, 1'd1} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd0, 5'd7, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd1, 5'd0, 1'd1} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd1, 5'd1, 1'd1} : icp_lc_expected = 5'b01101;
  {SERDES, 4'd1, 5'd2, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd1, 5'd3, 1'd1} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd1, 5'd4, 1'd1} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd1, 5'd5, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd1, 5'd6, 1'd1} : icp_lc_expected = 5'b00111;
  {SERDES, 4'd1, 5'd7, 1'd1} : icp_lc_expected = 5'b00110;
  {SERDES, 4'd2, 5'd0, 1'd1} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd2, 5'd1, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd2, 5'd2, 1'd1} : icp_lc_expected = 5'b01101;
  {SERDES, 4'd2, 5'd3, 1'd1} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd2, 5'd4, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd2, 5'd5, 1'd1} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd2, 5'd6, 1'd1} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd2, 5'd7, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd3, 5'd0, 1'd1} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd3, 5'd1, 1'd1} : icp_lc_expected = 5'b01101;
  {SERDES, 4'd3, 5'd2, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd3, 5'd3, 1'd1} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd3, 5'd4, 1'd1} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd3, 5'd5, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd3, 5'd6, 1'd1} : icp_lc_expected = 5'b00111;
  {SERDES, 4'd3, 5'd7, 1'd1} : icp_lc_expected = 5'b00110;
  {SERDES, 4'd4, 5'd0, 1'd1} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd4, 5'd1, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd4, 5'd2, 1'd1} : icp_lc_expected = 5'b01101;
  {SERDES, 4'd4, 5'd3, 1'd1} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd4, 5'd4, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd4, 5'd5, 1'd1} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd4, 5'd6, 1'd1} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd4, 5'd7, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd5, 5'd0, 1'd1} : icp_lc_expected = 5'b01101;
  {SERDES, 4'd5, 5'd1, 1'd1} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd5, 5'd2, 1'd1} : icp_lc_expected = 5'b01010;
  {SERDES, 4'd5, 5'd3, 1'd1} : icp_lc_expected = 5'b01101;
  {SERDES, 4'd5, 5'd4, 1'd1} : icp_lc_expected = 5'b01101;
  {SERDES, 4'd5, 5'd5, 1'd1} : icp_lc_expected = 5'b01010;
  {SERDES, 4'd5, 5'd6, 1'd1} : icp_lc_expected = 5'b01101;
  {SERDES, 4'd5, 5'd7, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd6, 5'd0, 1'd1} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd6, 5'd1, 1'd1} : icp_lc_expected = 5'b01101;
  {SERDES, 4'd6, 5'd2, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd6, 5'd3, 1'd1} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd6, 5'd4, 1'd1} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd6, 5'd5, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd6, 5'd6, 1'd1} : icp_lc_expected = 5'b00111;
  {SERDES, 4'd6, 5'd7, 1'd1} : icp_lc_expected = 5'b00110;
  {SERDES, 4'd7, 5'd0, 1'd1} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd7, 5'd1, 1'd1} : icp_lc_expected = 5'b01101;
  {SERDES, 4'd7, 5'd2, 1'd1} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd7, 5'd3, 1'd1} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd7, 5'd4, 1'd1} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd7, 5'd5, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd7, 5'd6, 1'd1} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd7, 5'd7, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd8, 5'd0, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd8, 5'd1, 1'd1} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd8, 5'd2, 1'd1} : icp_lc_expected = 5'b01010;
  {SERDES, 4'd8, 5'd3, 1'd1} : icp_lc_expected = 5'b01001;
  {SERDES, 4'd8, 5'd4, 1'd1} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd8, 5'd5, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd8, 5'd6, 1'd1} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd8, 5'd7, 1'd1} : icp_lc_expected = 5'b01001;
  {SERDES, 4'd9, 5'd0, 1'd1} : icp_lc_expected = 5'b01101;
  {SERDES, 4'd9, 5'd1, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd9, 5'd2, 1'd1} : icp_lc_expected = 5'b01011;
  {SERDES, 4'd9, 5'd3, 1'd1} : icp_lc_expected = 5'b01001;
  {SERDES, 4'd9, 5'd4, 1'd1} : icp_lc_expected = 5'b01010;
  {SERDES, 4'd9, 5'd5, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd9, 5'd6, 1'd1} : icp_lc_expected = 5'b01010;
  {SERDES, 4'd9, 5'd7, 1'd1} : icp_lc_expected = 5'b01001;
  {SERDES, 4'd12, 5'd0, 1'd1} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd12, 5'd1, 1'd1} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd12, 5'd2, 1'd1} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd12, 5'd3, 1'd1} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd12, 5'd4, 1'd1} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd12, 5'd5, 1'd1} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd12, 5'd6, 1'd1} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd12, 5'd7, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd13, 5'd0, 1'd1} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd13, 5'd1, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd13, 5'd2, 1'd1} : icp_lc_expected = 5'b01101;
  {SERDES, 4'd13, 5'd3, 1'd1} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd13, 5'd4, 1'd1} : icp_lc_expected = 5'b01100;
  {SERDES, 4'd13, 5'd5, 1'd1} : icp_lc_expected = 5'b01110;
  {SERDES, 4'd13, 5'd6, 1'd1} : icp_lc_expected = 5'b01111;
  {SERDES, 4'd13, 5'd7, 1'd1} : icp_lc_expected = 5'b01100;
  {SAS, 4'd0, 5'd0, 1'd1} : icp_lc_expected = 5'b01111;
  {SAS, 4'd0, 5'd1, 1'd1} : icp_lc_expected = 5'b01111;
  {SAS, 4'd0, 5'd2, 1'd1} : icp_lc_expected = 5'b01000;
  {SAS, 4'd0, 5'd3, 1'd1} : icp_lc_expected = 5'b01010;
  {SAS, 4'd0, 5'd4, 1'd1} : icp_lc_expected = 5'b01010;
  {SAS, 4'd0, 5'd5, 1'd1} : icp_lc_expected = 5'b01100;
  {SAS, 4'd0, 5'd6, 1'd1} : icp_lc_expected = 5'b01001;
  {SAS, 4'd0, 5'd7, 1'd1} : icp_lc_expected = 5'b01101;
  {SAS, 4'd1, 5'd0, 1'd1} : icp_lc_expected = 5'b01111;
  {SAS, 4'd1, 5'd1, 1'd1} : icp_lc_expected = 5'b01111;
  {SAS, 4'd1, 5'd2, 1'd1} : icp_lc_expected = 5'b01000;
  {SAS, 4'd1, 5'd3, 1'd1} : icp_lc_expected = 5'b01010;
  {SAS, 4'd1, 5'd4, 1'd1} : icp_lc_expected = 5'b01010;
  {SAS, 4'd1, 5'd5, 1'd1} : icp_lc_expected = 5'b01100;
  {SAS, 4'd1, 5'd6, 1'd1} : icp_lc_expected = 5'b01001;
  {SAS, 4'd1, 5'd7, 1'd1} : icp_lc_expected = 5'b01101;
  {SAS, 4'd2, 5'd0, 1'd1} : icp_lc_expected = 5'b01111;
  {SAS, 4'd2, 5'd1, 1'd1} : icp_lc_expected = 5'b01111;
  {SAS, 4'd2, 5'd2, 1'd1} : icp_lc_expected = 5'b01000;
  {SAS, 4'd2, 5'd3, 1'd1} : icp_lc_expected = 5'b01010;
  {SAS, 4'd2, 5'd4, 1'd1} : icp_lc_expected = 5'b01010;
  {SAS, 4'd2, 5'd5, 1'd1} : icp_lc_expected = 5'b01100;
  {SAS, 4'd2, 5'd6, 1'd1} : icp_lc_expected = 5'b01001;
  {SAS, 4'd2, 5'd7, 1'd1} : icp_lc_expected = 5'b01101;
  {SAS, 4'd3, 5'd0, 1'd1} : icp_lc_expected = 5'b01111;
  {SAS, 4'd3, 5'd1, 1'd1} : icp_lc_expected = 5'b01111;
  {SAS, 4'd3, 5'd2, 1'd1} : icp_lc_expected = 5'b01000;
  {SAS, 4'd3, 5'd3, 1'd1} : icp_lc_expected = 5'b01010;
  {SAS, 4'd3, 5'd4, 1'd1} : icp_lc_expected = 5'b01010;
  {SAS, 4'd3, 5'd5, 1'd1} : icp_lc_expected = 5'b01100;
  {SAS, 4'd3, 5'd6, 1'd1} : icp_lc_expected = 5'b01001;
  {SAS, 4'd3, 5'd7, 1'd1} : icp_lc_expected = 5'b01101;
  {SAS, 4'd4, 5'd0, 1'd1} : icp_lc_expected = 5'b01111;
  {SAS, 4'd4, 5'd1, 1'd1} : icp_lc_expected = 5'b01111;
  {SAS, 4'd4, 5'd2, 1'd1} : icp_lc_expected = 5'b01101;
  {SAS, 4'd4, 5'd3, 1'd1} : icp_lc_expected = 5'b01100;
  {SAS, 4'd4, 5'd4, 1'd1} : icp_lc_expected = 5'b01110;
  {SAS, 4'd4, 5'd5, 1'd1} : icp_lc_expected = 5'b01100;
  {SAS, 4'd4, 5'd6, 1'd1} : icp_lc_expected = 5'b01101;
  {SAS, 4'd4, 5'd7, 1'd1} : icp_lc_expected = 5'b01100;
  {PCIE, 4'd2, 5'd0, 1'd1} : icp_lc_expected = 5'b01111;
  {PCIE, 4'd2, 5'd1, 1'd1} : icp_lc_expected = 5'b01110;
  {PCIE, 4'd2, 5'd2, 1'd1} : icp_lc_expected = 5'b01111;
  {PCIE, 4'd2, 5'd3, 1'd1} : icp_lc_expected = 5'b01111;
  {PCIE, 4'd2, 5'd4, 1'd1} : icp_lc_expected = 5'b01101;
  {PCIE, 4'd2, 5'd5, 1'd1} : icp_lc_expected = 5'b01111;
  {PCIE, 4'd2, 5'd6, 1'd1} : icp_lc_expected = 5'b01011;
  {PCIE, 4'd2, 5'd7, 1'd1} : icp_lc_expected = 5'b01111;
  {PCIE, 4'd3, 5'd0, 1'd1} : icp_lc_expected = 5'b01111;
  {PCIE, 4'd3, 5'd1, 1'd1} : icp_lc_expected = 5'b01110;
  {PCIE, 4'd3, 5'd2, 1'd1} : icp_lc_expected = 5'b01111;
  {PCIE, 4'd3, 5'd3, 1'd1} : icp_lc_expected = 5'b01111;
  {PCIE, 4'd3, 5'd4, 1'd1} : icp_lc_expected = 5'b01101;
  {PCIE, 4'd3, 5'd5, 1'd1} : icp_lc_expected = 5'b01111;
  {PCIE, 4'd3, 5'd6, 1'd1} : icp_lc_expected = 5'b01011;
  {PCIE, 4'd3, 5'd7, 1'd1} : icp_lc_expected = 5'b01111;
default: icp_lc_expected = 5'bzzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel} )
  {USB, 4'd1, 5'd0, 1'd0} : pll_lpfr_expected = 2'b01;
  {USB, 4'd1, 5'd1, 1'd0} : pll_lpfr_expected = 2'b01;
  {USB, 4'd1, 5'd2, 1'd0} : pll_lpfr_expected = 2'b01;
  {USB, 4'd1, 5'd3, 1'd0} : pll_lpfr_expected = 2'b01;
  {USB, 4'd1, 5'd4, 1'd0} : pll_lpfr_expected = 2'b01;
  {USB, 4'd1, 5'd5, 1'd0} : pll_lpfr_expected = 2'b01;
  {USB, 4'd1, 5'd6, 1'd0} : pll_lpfr_expected = 2'b00;
  {USB, 4'd1, 5'd7, 1'd0} : pll_lpfr_expected = 2'b00;
  {USB, 4'd2, 5'd0, 1'd0} : pll_lpfr_expected = 2'b01;
  {USB, 4'd2, 5'd1, 1'd0} : pll_lpfr_expected = 2'b01;
  {USB, 4'd2, 5'd2, 1'd0} : pll_lpfr_expected = 2'b01;
  {USB, 4'd2, 5'd3, 1'd0} : pll_lpfr_expected = 2'b01;
  {USB, 4'd2, 5'd4, 1'd0} : pll_lpfr_expected = 2'b01;
  {USB, 4'd2, 5'd5, 1'd0} : pll_lpfr_expected = 2'b01;
  {USB, 4'd2, 5'd6, 1'd0} : pll_lpfr_expected = 2'b00;
  {USB, 4'd2, 5'd7, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd0, 5'd0, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd0, 5'd1, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd0, 5'd2, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd0, 5'd3, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd0, 5'd4, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd0, 5'd5, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd0, 5'd6, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd0, 5'd7, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd1, 5'd0, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd1, 5'd1, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd1, 5'd2, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd1, 5'd3, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd1, 5'd4, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd1, 5'd5, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd1, 5'd6, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd1, 5'd7, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd2, 5'd0, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd2, 5'd1, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd2, 5'd2, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd2, 5'd3, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd2, 5'd4, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd2, 5'd5, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd2, 5'd6, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd2, 5'd7, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd3, 5'd0, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd3, 5'd1, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd3, 5'd2, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd3, 5'd3, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd3, 5'd4, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd3, 5'd5, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd3, 5'd6, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd3, 5'd7, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd4, 5'd0, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd4, 5'd1, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd4, 5'd2, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd4, 5'd3, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd4, 5'd4, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd4, 5'd5, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd4, 5'd6, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd4, 5'd7, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd5, 5'd0, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd5, 5'd1, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd5, 5'd2, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd5, 5'd3, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd5, 5'd4, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd5, 5'd5, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd5, 5'd6, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd5, 5'd7, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd6, 5'd0, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd6, 5'd1, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd6, 5'd2, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd6, 5'd3, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd6, 5'd4, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd6, 5'd5, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd6, 5'd6, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd6, 5'd7, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd7, 5'd0, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd7, 5'd1, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd7, 5'd2, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd7, 5'd3, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd7, 5'd4, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd7, 5'd5, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd7, 5'd6, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd7, 5'd7, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd8, 5'd0, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd8, 5'd1, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd8, 5'd2, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd8, 5'd3, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd8, 5'd4, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd8, 5'd5, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd8, 5'd6, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd8, 5'd7, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd9, 5'd0, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd9, 5'd1, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd9, 5'd2, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd9, 5'd3, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd9, 5'd4, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd9, 5'd5, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd9, 5'd6, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd9, 5'd7, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd12, 5'd0, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd12, 5'd1, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd12, 5'd2, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd12, 5'd3, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd12, 5'd4, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd12, 5'd5, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd12, 5'd6, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd12, 5'd7, 1'd0} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd13, 5'd0, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd13, 5'd1, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd13, 5'd2, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd13, 5'd3, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd13, 5'd4, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd13, 5'd5, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd13, 5'd6, 1'd0} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd13, 5'd7, 1'd0} : pll_lpfr_expected = 2'b00;
  {SAS, 4'd0, 5'd0, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd0, 5'd1, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd0, 5'd2, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd0, 5'd3, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd0, 5'd4, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd0, 5'd5, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd0, 5'd6, 1'd0} : pll_lpfr_expected = 2'b00;
  {SAS, 4'd0, 5'd7, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd1, 5'd0, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd1, 5'd1, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd1, 5'd2, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd1, 5'd3, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd1, 5'd4, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd1, 5'd5, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd1, 5'd6, 1'd0} : pll_lpfr_expected = 2'b00;
  {SAS, 4'd1, 5'd7, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd2, 5'd0, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd2, 5'd1, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd2, 5'd2, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd2, 5'd3, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd2, 5'd4, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd2, 5'd5, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd2, 5'd6, 1'd0} : pll_lpfr_expected = 2'b00;
  {SAS, 4'd2, 5'd7, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd3, 5'd0, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd3, 5'd1, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd3, 5'd2, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd3, 5'd3, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd3, 5'd4, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd3, 5'd5, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd3, 5'd6, 1'd0} : pll_lpfr_expected = 2'b00;
  {SAS, 4'd3, 5'd7, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd4, 5'd0, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd4, 5'd1, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd4, 5'd2, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd4, 5'd3, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd4, 5'd4, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd4, 5'd5, 1'd0} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd4, 5'd6, 1'd0} : pll_lpfr_expected = 2'b00;
  {SAS, 4'd4, 5'd7, 1'd0} : pll_lpfr_expected = 2'b00;
  {PCIE, 4'd2, 5'd0, 1'd0} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd2, 5'd1, 1'd0} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd2, 5'd2, 1'd0} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd2, 5'd3, 1'd0} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd2, 5'd4, 1'd0} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd2, 5'd5, 1'd0} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd2, 5'd6, 1'd0} : pll_lpfr_expected = 2'b00;
  {PCIE, 4'd2, 5'd7, 1'd0} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd3, 5'd0, 1'd0} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd3, 5'd1, 1'd0} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd3, 5'd2, 1'd0} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd3, 5'd3, 1'd0} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd3, 5'd4, 1'd0} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd3, 5'd5, 1'd0} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd3, 5'd6, 1'd0} : pll_lpfr_expected = 2'b00;
  {PCIE, 4'd3, 5'd7, 1'd0} : pll_lpfr_expected = 2'b01;
  {USB, 4'd1, 5'd0, 1'd1} : pll_lpfr_expected = 2'b01;
  {USB, 4'd1, 5'd1, 1'd1} : pll_lpfr_expected = 2'b01;
  {USB, 4'd1, 5'd2, 1'd1} : pll_lpfr_expected = 2'b01;
  {USB, 4'd1, 5'd3, 1'd1} : pll_lpfr_expected = 2'b01;
  {USB, 4'd1, 5'd4, 1'd1} : pll_lpfr_expected = 2'b01;
  {USB, 4'd1, 5'd5, 1'd1} : pll_lpfr_expected = 2'b01;
  {USB, 4'd1, 5'd6, 1'd1} : pll_lpfr_expected = 2'b00;
  {USB, 4'd1, 5'd7, 1'd1} : pll_lpfr_expected = 2'b00;
  {USB, 4'd2, 5'd0, 1'd1} : pll_lpfr_expected = 2'b01;
  {USB, 4'd2, 5'd1, 1'd1} : pll_lpfr_expected = 2'b01;
  {USB, 4'd2, 5'd2, 1'd1} : pll_lpfr_expected = 2'b01;
  {USB, 4'd2, 5'd3, 1'd1} : pll_lpfr_expected = 2'b01;
  {USB, 4'd2, 5'd4, 1'd1} : pll_lpfr_expected = 2'b01;
  {USB, 4'd2, 5'd5, 1'd1} : pll_lpfr_expected = 2'b01;
  {USB, 4'd2, 5'd6, 1'd1} : pll_lpfr_expected = 2'b00;
  {USB, 4'd2, 5'd7, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd0, 5'd0, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd0, 5'd1, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd0, 5'd2, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd0, 5'd3, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd0, 5'd4, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd0, 5'd5, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd0, 5'd6, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd0, 5'd7, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd1, 5'd0, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd1, 5'd1, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd1, 5'd2, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd1, 5'd3, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd1, 5'd4, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd1, 5'd5, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd1, 5'd6, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd1, 5'd7, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd2, 5'd0, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd2, 5'd1, 1'd1} : pll_lpfr_expected = 2'b10;
  {SERDES, 4'd2, 5'd2, 1'd1} : pll_lpfr_expected = 2'b10;
  {SERDES, 4'd2, 5'd3, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd2, 5'd4, 1'd1} : pll_lpfr_expected = 2'b10;
  {SERDES, 4'd2, 5'd5, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd2, 5'd6, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd2, 5'd7, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd3, 5'd0, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd3, 5'd1, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd3, 5'd2, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd3, 5'd3, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd3, 5'd4, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd3, 5'd5, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd3, 5'd6, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd3, 5'd7, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd4, 5'd0, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd4, 5'd1, 1'd1} : pll_lpfr_expected = 2'b10;
  {SERDES, 4'd4, 5'd2, 1'd1} : pll_lpfr_expected = 2'b10;
  {SERDES, 4'd4, 5'd3, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd4, 5'd4, 1'd1} : pll_lpfr_expected = 2'b10;
  {SERDES, 4'd4, 5'd5, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd4, 5'd6, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd4, 5'd7, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd5, 5'd0, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd5, 5'd1, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd5, 5'd2, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd5, 5'd3, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd5, 5'd4, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd5, 5'd5, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd5, 5'd6, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd5, 5'd7, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd6, 5'd0, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd6, 5'd1, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd6, 5'd2, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd6, 5'd3, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd6, 5'd4, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd6, 5'd5, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd6, 5'd6, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd6, 5'd7, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd7, 5'd0, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd7, 5'd1, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd7, 5'd2, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd7, 5'd3, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd7, 5'd4, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd7, 5'd5, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd7, 5'd6, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd7, 5'd7, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd8, 5'd0, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd8, 5'd1, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd8, 5'd2, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd8, 5'd3, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd8, 5'd4, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd8, 5'd5, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd8, 5'd6, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd8, 5'd7, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd9, 5'd0, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd9, 5'd1, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd9, 5'd2, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd9, 5'd3, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd9, 5'd4, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd9, 5'd5, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd9, 5'd6, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd9, 5'd7, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd12, 5'd0, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd12, 5'd1, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd12, 5'd2, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd12, 5'd3, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd12, 5'd4, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd12, 5'd5, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd12, 5'd6, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd12, 5'd7, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd13, 5'd0, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd13, 5'd1, 1'd1} : pll_lpfr_expected = 2'b10;
  {SERDES, 4'd13, 5'd2, 1'd1} : pll_lpfr_expected = 2'b10;
  {SERDES, 4'd13, 5'd3, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd13, 5'd4, 1'd1} : pll_lpfr_expected = 2'b10;
  {SERDES, 4'd13, 5'd5, 1'd1} : pll_lpfr_expected = 2'b01;
  {SERDES, 4'd13, 5'd6, 1'd1} : pll_lpfr_expected = 2'b00;
  {SERDES, 4'd13, 5'd7, 1'd1} : pll_lpfr_expected = 2'b00;
  {SAS, 4'd0, 5'd0, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd0, 5'd1, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd0, 5'd2, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd0, 5'd3, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd0, 5'd4, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd0, 5'd5, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd0, 5'd6, 1'd1} : pll_lpfr_expected = 2'b00;
  {SAS, 4'd0, 5'd7, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd1, 5'd0, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd1, 5'd1, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd1, 5'd2, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd1, 5'd3, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd1, 5'd4, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd1, 5'd5, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd1, 5'd6, 1'd1} : pll_lpfr_expected = 2'b00;
  {SAS, 4'd1, 5'd7, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd2, 5'd0, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd2, 5'd1, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd2, 5'd2, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd2, 5'd3, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd2, 5'd4, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd2, 5'd5, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd2, 5'd6, 1'd1} : pll_lpfr_expected = 2'b00;
  {SAS, 4'd2, 5'd7, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd3, 5'd0, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd3, 5'd1, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd3, 5'd2, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd3, 5'd3, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd3, 5'd4, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd3, 5'd5, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd3, 5'd6, 1'd1} : pll_lpfr_expected = 2'b00;
  {SAS, 4'd3, 5'd7, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd4, 5'd0, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd4, 5'd1, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd4, 5'd2, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd4, 5'd3, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd4, 5'd4, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd4, 5'd5, 1'd1} : pll_lpfr_expected = 2'b01;
  {SAS, 4'd4, 5'd6, 1'd1} : pll_lpfr_expected = 2'b00;
  {SAS, 4'd4, 5'd7, 1'd1} : pll_lpfr_expected = 2'b00;
  {PCIE, 4'd2, 5'd0, 1'd1} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd2, 5'd1, 1'd1} : pll_lpfr_expected = 2'b10;
  {PCIE, 4'd2, 5'd2, 1'd1} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd2, 5'd3, 1'd1} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd2, 5'd4, 1'd1} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd2, 5'd5, 1'd1} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd2, 5'd6, 1'd1} : pll_lpfr_expected = 2'b00;
  {PCIE, 4'd2, 5'd7, 1'd1} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd3, 5'd0, 1'd1} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd3, 5'd1, 1'd1} : pll_lpfr_expected = 2'b10;
  {PCIE, 4'd3, 5'd2, 1'd1} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd3, 5'd3, 1'd1} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd3, 5'd4, 1'd1} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd3, 5'd5, 1'd1} : pll_lpfr_expected = 2'b01;
  {PCIE, 4'd3, 5'd6, 1'd1} : pll_lpfr_expected = 2'b00;
  {PCIE, 4'd3, 5'd7, 1'd1} : pll_lpfr_expected = 2'b01;
default: pll_lpfr_expected = 2'bzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel} )
  {USB, 4'd1, 5'd0, 1'd0} : pll_lpfc_expected = 2'b01;
  {USB, 4'd1, 5'd1, 1'd0} : pll_lpfc_expected = 2'b01;
  {USB, 4'd1, 5'd2, 1'd0} : pll_lpfc_expected = 2'b01;
  {USB, 4'd1, 5'd3, 1'd0} : pll_lpfc_expected = 2'b01;
  {USB, 4'd1, 5'd4, 1'd0} : pll_lpfc_expected = 2'b01;
  {USB, 4'd1, 5'd5, 1'd0} : pll_lpfc_expected = 2'b01;
  {USB, 4'd1, 5'd6, 1'd0} : pll_lpfc_expected = 2'b01;
  {USB, 4'd1, 5'd7, 1'd0} : pll_lpfc_expected = 2'b01;
  {USB, 4'd2, 5'd0, 1'd0} : pll_lpfc_expected = 2'b01;
  {USB, 4'd2, 5'd1, 1'd0} : pll_lpfc_expected = 2'b01;
  {USB, 4'd2, 5'd2, 1'd0} : pll_lpfc_expected = 2'b01;
  {USB, 4'd2, 5'd3, 1'd0} : pll_lpfc_expected = 2'b01;
  {USB, 4'd2, 5'd4, 1'd0} : pll_lpfc_expected = 2'b01;
  {USB, 4'd2, 5'd5, 1'd0} : pll_lpfc_expected = 2'b01;
  {USB, 4'd2, 5'd6, 1'd0} : pll_lpfc_expected = 2'b01;
  {USB, 4'd2, 5'd7, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd0, 5'd0, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd0, 5'd1, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd0, 5'd2, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd0, 5'd3, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd0, 5'd4, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd0, 5'd5, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd0, 5'd6, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd0, 5'd7, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd1, 5'd0, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd1, 5'd1, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd1, 5'd2, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd1, 5'd3, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd1, 5'd4, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd1, 5'd5, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd1, 5'd6, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd1, 5'd7, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd2, 5'd0, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd2, 5'd1, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd2, 5'd2, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd2, 5'd3, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd2, 5'd4, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd2, 5'd5, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd2, 5'd6, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd2, 5'd7, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd3, 5'd0, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd3, 5'd1, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd3, 5'd2, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd3, 5'd3, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd3, 5'd4, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd3, 5'd5, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd3, 5'd6, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd3, 5'd7, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd4, 5'd0, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd4, 5'd1, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd4, 5'd2, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd4, 5'd3, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd4, 5'd4, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd4, 5'd5, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd4, 5'd6, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd4, 5'd7, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd5, 5'd0, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd5, 5'd1, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd5, 5'd2, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd5, 5'd3, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd5, 5'd4, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd5, 5'd5, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd5, 5'd6, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd5, 5'd7, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd6, 5'd0, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd6, 5'd1, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd6, 5'd2, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd6, 5'd3, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd6, 5'd4, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd6, 5'd5, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd6, 5'd6, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd6, 5'd7, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd7, 5'd0, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd7, 5'd1, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd7, 5'd2, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd7, 5'd3, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd7, 5'd4, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd7, 5'd5, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd7, 5'd6, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd7, 5'd7, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd8, 5'd0, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd8, 5'd1, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd8, 5'd2, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd8, 5'd3, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd8, 5'd4, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd8, 5'd5, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd8, 5'd6, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd8, 5'd7, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd9, 5'd0, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd9, 5'd1, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd9, 5'd2, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd9, 5'd3, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd9, 5'd4, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd9, 5'd5, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd9, 5'd6, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd9, 5'd7, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd12, 5'd0, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd12, 5'd1, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd12, 5'd2, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd12, 5'd3, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd12, 5'd4, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd12, 5'd5, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd12, 5'd6, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd12, 5'd7, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd13, 5'd0, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd13, 5'd1, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd13, 5'd2, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd13, 5'd3, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd13, 5'd4, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd13, 5'd5, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd13, 5'd6, 1'd0} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd13, 5'd7, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd0, 5'd0, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd0, 5'd1, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd0, 5'd2, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd0, 5'd3, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd0, 5'd4, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd0, 5'd5, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd0, 5'd6, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd0, 5'd7, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd1, 5'd0, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd1, 5'd1, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd1, 5'd2, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd1, 5'd3, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd1, 5'd4, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd1, 5'd5, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd1, 5'd6, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd1, 5'd7, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd2, 5'd0, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd2, 5'd1, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd2, 5'd2, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd2, 5'd3, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd2, 5'd4, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd2, 5'd5, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd2, 5'd6, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd2, 5'd7, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd3, 5'd0, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd3, 5'd1, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd3, 5'd2, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd3, 5'd3, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd3, 5'd4, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd3, 5'd5, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd3, 5'd6, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd3, 5'd7, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd4, 5'd0, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd4, 5'd1, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd4, 5'd2, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd4, 5'd3, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd4, 5'd4, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd4, 5'd5, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd4, 5'd6, 1'd0} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd4, 5'd7, 1'd0} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd2, 5'd0, 1'd0} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd2, 5'd1, 1'd0} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd2, 5'd2, 1'd0} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd2, 5'd3, 1'd0} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd2, 5'd4, 1'd0} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd2, 5'd5, 1'd0} : pll_lpfc_expected = 2'b00;
  {PCIE, 4'd2, 5'd6, 1'd0} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd2, 5'd7, 1'd0} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd3, 5'd0, 1'd0} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd3, 5'd1, 1'd0} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd3, 5'd2, 1'd0} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd3, 5'd3, 1'd0} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd3, 5'd4, 1'd0} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd3, 5'd5, 1'd0} : pll_lpfc_expected = 2'b00;
  {PCIE, 4'd3, 5'd6, 1'd0} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd3, 5'd7, 1'd0} : pll_lpfc_expected = 2'b01;
  {USB, 4'd1, 5'd0, 1'd1} : pll_lpfc_expected = 2'b01;
  {USB, 4'd1, 5'd1, 1'd1} : pll_lpfc_expected = 2'b01;
  {USB, 4'd1, 5'd2, 1'd1} : pll_lpfc_expected = 2'b01;
  {USB, 4'd1, 5'd3, 1'd1} : pll_lpfc_expected = 2'b01;
  {USB, 4'd1, 5'd4, 1'd1} : pll_lpfc_expected = 2'b01;
  {USB, 4'd1, 5'd5, 1'd1} : pll_lpfc_expected = 2'b01;
  {USB, 4'd1, 5'd6, 1'd1} : pll_lpfc_expected = 2'b01;
  {USB, 4'd1, 5'd7, 1'd1} : pll_lpfc_expected = 2'b01;
  {USB, 4'd2, 5'd0, 1'd1} : pll_lpfc_expected = 2'b01;
  {USB, 4'd2, 5'd1, 1'd1} : pll_lpfc_expected = 2'b01;
  {USB, 4'd2, 5'd2, 1'd1} : pll_lpfc_expected = 2'b01;
  {USB, 4'd2, 5'd3, 1'd1} : pll_lpfc_expected = 2'b01;
  {USB, 4'd2, 5'd4, 1'd1} : pll_lpfc_expected = 2'b01;
  {USB, 4'd2, 5'd5, 1'd1} : pll_lpfc_expected = 2'b01;
  {USB, 4'd2, 5'd6, 1'd1} : pll_lpfc_expected = 2'b01;
  {USB, 4'd2, 5'd7, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd0, 5'd0, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd0, 5'd1, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd0, 5'd2, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd0, 5'd3, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd0, 5'd4, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd0, 5'd5, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd0, 5'd6, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd0, 5'd7, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd1, 5'd0, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd1, 5'd1, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd1, 5'd2, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd1, 5'd3, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd1, 5'd4, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd1, 5'd5, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd1, 5'd6, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd1, 5'd7, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd2, 5'd0, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd2, 5'd1, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd2, 5'd2, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd2, 5'd3, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd2, 5'd4, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd2, 5'd5, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd2, 5'd6, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd2, 5'd7, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd3, 5'd0, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd3, 5'd1, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd3, 5'd2, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd3, 5'd3, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd3, 5'd4, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd3, 5'd5, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd3, 5'd6, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd3, 5'd7, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd4, 5'd0, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd4, 5'd1, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd4, 5'd2, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd4, 5'd3, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd4, 5'd4, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd4, 5'd5, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd4, 5'd6, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd4, 5'd7, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd5, 5'd0, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd5, 5'd1, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd5, 5'd2, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd5, 5'd3, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd5, 5'd4, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd5, 5'd5, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd5, 5'd6, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd5, 5'd7, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd6, 5'd0, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd6, 5'd1, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd6, 5'd2, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd6, 5'd3, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd6, 5'd4, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd6, 5'd5, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd6, 5'd6, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd6, 5'd7, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd7, 5'd0, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd7, 5'd1, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd7, 5'd2, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd7, 5'd3, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd7, 5'd4, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd7, 5'd5, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd7, 5'd6, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd7, 5'd7, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd8, 5'd0, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd8, 5'd1, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd8, 5'd2, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd8, 5'd3, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd8, 5'd4, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd8, 5'd5, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd8, 5'd6, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd8, 5'd7, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd9, 5'd0, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd9, 5'd1, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd9, 5'd2, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd9, 5'd3, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd9, 5'd4, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd9, 5'd5, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd9, 5'd6, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd9, 5'd7, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd12, 5'd0, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd12, 5'd1, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd12, 5'd2, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd12, 5'd3, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd12, 5'd4, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd12, 5'd5, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd12, 5'd6, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd12, 5'd7, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd13, 5'd0, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd13, 5'd1, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd13, 5'd2, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd13, 5'd3, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd13, 5'd4, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd13, 5'd5, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd13, 5'd6, 1'd1} : pll_lpfc_expected = 2'b01;
  {SERDES, 4'd13, 5'd7, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd0, 5'd0, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd0, 5'd1, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd0, 5'd2, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd0, 5'd3, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd0, 5'd4, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd0, 5'd5, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd0, 5'd6, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd0, 5'd7, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd1, 5'd0, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd1, 5'd1, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd1, 5'd2, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd1, 5'd3, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd1, 5'd4, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd1, 5'd5, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd1, 5'd6, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd1, 5'd7, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd2, 5'd0, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd2, 5'd1, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd2, 5'd2, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd2, 5'd3, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd2, 5'd4, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd2, 5'd5, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd2, 5'd6, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd2, 5'd7, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd3, 5'd0, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd3, 5'd1, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd3, 5'd2, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd3, 5'd3, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd3, 5'd4, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd3, 5'd5, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd3, 5'd6, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd3, 5'd7, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd4, 5'd0, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd4, 5'd1, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd4, 5'd2, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd4, 5'd3, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd4, 5'd4, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd4, 5'd5, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd4, 5'd6, 1'd1} : pll_lpfc_expected = 2'b01;
  {SAS, 4'd4, 5'd7, 1'd1} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd2, 5'd0, 1'd1} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd2, 5'd1, 1'd1} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd2, 5'd2, 1'd1} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd2, 5'd3, 1'd1} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd2, 5'd4, 1'd1} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd2, 5'd5, 1'd1} : pll_lpfc_expected = 2'b00;
  {PCIE, 4'd2, 5'd6, 1'd1} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd2, 5'd7, 1'd1} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd3, 5'd0, 1'd1} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd3, 5'd1, 1'd1} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd3, 5'd2, 1'd1} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd3, 5'd3, 1'd1} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd3, 5'd4, 1'd1} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd3, 5'd5, 1'd1} : pll_lpfc_expected = 2'b00;
  {PCIE, 4'd3, 5'd6, 1'd1} : pll_lpfc_expected = 2'b01;
  {PCIE, 4'd3, 5'd7, 1'd1} : pll_lpfc_expected = 2'b01;
default: pll_lpfc_expected = 2'bzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel} )
  {USB, 4'd1, 5'd0, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd1, 5'd1, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd1, 5'd2, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd1, 5'd3, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd1, 5'd4, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd1, 5'd5, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd1, 5'd6, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd1, 5'd7, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd2, 5'd0, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd2, 5'd1, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd2, 5'd2, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd2, 5'd3, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd2, 5'd4, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd2, 5'd5, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd2, 5'd6, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd2, 5'd7, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd0, 5'd0, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd0, 5'd1, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd0, 5'd2, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd0, 5'd3, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd0, 5'd4, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd0, 5'd5, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd0, 5'd6, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd0, 5'd7, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd1, 5'd0, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd1, 5'd1, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd1, 5'd2, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd1, 5'd3, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd1, 5'd4, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd1, 5'd5, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd1, 5'd6, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd1, 5'd7, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd2, 5'd0, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd2, 5'd1, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd2, 5'd2, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd2, 5'd3, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd2, 5'd4, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd2, 5'd5, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd2, 5'd6, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd2, 5'd7, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd3, 5'd0, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd3, 5'd1, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd3, 5'd2, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd3, 5'd3, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd3, 5'd4, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd3, 5'd5, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd3, 5'd6, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd3, 5'd7, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd4, 5'd0, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd4, 5'd1, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd4, 5'd2, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd4, 5'd3, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd4, 5'd4, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd4, 5'd5, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd4, 5'd6, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd4, 5'd7, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd5, 5'd0, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd5, 5'd1, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd5, 5'd2, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd5, 5'd3, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd5, 5'd4, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd5, 5'd5, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd5, 5'd6, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd5, 5'd7, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd6, 5'd0, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd6, 5'd1, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd6, 5'd2, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd6, 5'd3, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd6, 5'd4, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd6, 5'd5, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd6, 5'd6, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd6, 5'd7, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd7, 5'd0, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd7, 5'd1, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd7, 5'd2, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd7, 5'd3, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd7, 5'd4, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd7, 5'd5, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd7, 5'd6, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd7, 5'd7, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd8, 5'd0, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd8, 5'd1, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd8, 5'd2, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd8, 5'd3, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd8, 5'd4, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd8, 5'd5, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd8, 5'd6, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd8, 5'd7, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd9, 5'd0, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd9, 5'd1, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd9, 5'd2, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd9, 5'd3, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd9, 5'd4, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd9, 5'd5, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd9, 5'd6, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd9, 5'd7, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd12, 5'd0, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd12, 5'd1, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd12, 5'd2, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd12, 5'd3, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd12, 5'd4, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd12, 5'd5, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd12, 5'd6, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd12, 5'd7, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd13, 5'd0, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd13, 5'd1, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd13, 5'd2, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd13, 5'd3, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd13, 5'd4, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd13, 5'd5, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd13, 5'd6, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd13, 5'd7, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SAS, 4'd0, 5'd0, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd0, 5'd1, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd0, 5'd2, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd0, 5'd3, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd0, 5'd4, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd0, 5'd5, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd0, 5'd6, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd0, 5'd7, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd1, 5'd0, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd1, 5'd1, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd1, 5'd2, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd1, 5'd3, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd1, 5'd4, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd1, 5'd5, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd1, 5'd6, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd1, 5'd7, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd2, 5'd0, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd2, 5'd1, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd2, 5'd2, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd2, 5'd3, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd2, 5'd4, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd2, 5'd5, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd2, 5'd6, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd2, 5'd7, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd3, 5'd0, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd3, 5'd1, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd3, 5'd2, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd3, 5'd3, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd3, 5'd4, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd3, 5'd5, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd3, 5'd6, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd3, 5'd7, 1'd0} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd4, 5'd0, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SAS, 4'd4, 5'd1, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SAS, 4'd4, 5'd2, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SAS, 4'd4, 5'd3, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SAS, 4'd4, 5'd4, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SAS, 4'd4, 5'd5, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SAS, 4'd4, 5'd6, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {SAS, 4'd4, 5'd7, 1'd0} : intpi_lcpll_expected = 4'b0100;
  {PCIE, 4'd2, 5'd0, 1'd0} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd2, 5'd1, 1'd0} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd2, 5'd2, 1'd0} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd2, 5'd3, 1'd0} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd2, 5'd4, 1'd0} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd2, 5'd5, 1'd0} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd2, 5'd6, 1'd0} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd2, 5'd7, 1'd0} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd3, 5'd0, 1'd0} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd3, 5'd1, 1'd0} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd3, 5'd2, 1'd0} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd3, 5'd3, 1'd0} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd3, 5'd4, 1'd0} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd3, 5'd5, 1'd0} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd3, 5'd6, 1'd0} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd3, 5'd7, 1'd0} : intpi_lcpll_expected = 4'b0011;
  {USB, 4'd1, 5'd0, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd1, 5'd1, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd1, 5'd2, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd1, 5'd3, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd1, 5'd4, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd1, 5'd5, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd1, 5'd6, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd1, 5'd7, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd2, 5'd0, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd2, 5'd1, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd2, 5'd2, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd2, 5'd3, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd2, 5'd4, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd2, 5'd5, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd2, 5'd6, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {USB, 4'd2, 5'd7, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd0, 5'd0, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd0, 5'd1, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd0, 5'd2, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd0, 5'd3, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd0, 5'd4, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd0, 5'd5, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd0, 5'd6, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd0, 5'd7, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd1, 5'd0, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd1, 5'd1, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd1, 5'd2, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd1, 5'd3, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd1, 5'd4, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd1, 5'd5, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd1, 5'd6, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd1, 5'd7, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd2, 5'd0, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd2, 5'd1, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd2, 5'd2, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd2, 5'd3, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd2, 5'd4, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd2, 5'd5, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd2, 5'd6, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd2, 5'd7, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd3, 5'd0, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd3, 5'd1, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd3, 5'd2, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd3, 5'd3, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd3, 5'd4, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd3, 5'd5, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd3, 5'd6, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd3, 5'd7, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd4, 5'd0, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd4, 5'd1, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd4, 5'd2, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd4, 5'd3, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd4, 5'd4, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd4, 5'd5, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd4, 5'd6, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd4, 5'd7, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd5, 5'd0, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd5, 5'd1, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd5, 5'd2, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd5, 5'd3, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd5, 5'd4, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd5, 5'd5, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd5, 5'd6, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd5, 5'd7, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd6, 5'd0, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd6, 5'd1, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd6, 5'd2, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd6, 5'd3, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd6, 5'd4, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd6, 5'd5, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd6, 5'd6, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd6, 5'd7, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd7, 5'd0, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd7, 5'd1, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd7, 5'd2, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd7, 5'd3, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd7, 5'd4, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd7, 5'd5, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd7, 5'd6, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd7, 5'd7, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd8, 5'd0, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd8, 5'd1, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd8, 5'd2, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd8, 5'd3, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd8, 5'd4, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd8, 5'd5, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd8, 5'd6, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd8, 5'd7, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd9, 5'd0, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd9, 5'd1, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd9, 5'd2, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd9, 5'd3, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd9, 5'd4, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd9, 5'd5, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd9, 5'd6, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd9, 5'd7, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SERDES, 4'd12, 5'd0, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd12, 5'd1, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd12, 5'd2, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd12, 5'd3, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd12, 5'd4, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd12, 5'd5, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd12, 5'd6, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd12, 5'd7, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd13, 5'd0, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd13, 5'd1, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd13, 5'd2, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd13, 5'd3, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd13, 5'd4, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd13, 5'd5, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd13, 5'd6, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SERDES, 4'd13, 5'd7, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SAS, 4'd0, 5'd0, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd0, 5'd1, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd0, 5'd2, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd0, 5'd3, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd0, 5'd4, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd0, 5'd5, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd0, 5'd6, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd0, 5'd7, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd1, 5'd0, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd1, 5'd1, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd1, 5'd2, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd1, 5'd3, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd1, 5'd4, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd1, 5'd5, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd1, 5'd6, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd1, 5'd7, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd2, 5'd0, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd2, 5'd1, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd2, 5'd2, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd2, 5'd3, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd2, 5'd4, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd2, 5'd5, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd2, 5'd6, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd2, 5'd7, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd3, 5'd0, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd3, 5'd1, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd3, 5'd2, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd3, 5'd3, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd3, 5'd4, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd3, 5'd5, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd3, 5'd6, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd3, 5'd7, 1'd1} : intpi_lcpll_expected = 4'b0110;
  {SAS, 4'd4, 5'd0, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SAS, 4'd4, 5'd1, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SAS, 4'd4, 5'd2, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SAS, 4'd4, 5'd3, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SAS, 4'd4, 5'd4, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SAS, 4'd4, 5'd5, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SAS, 4'd4, 5'd6, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {SAS, 4'd4, 5'd7, 1'd1} : intpi_lcpll_expected = 4'b0100;
  {PCIE, 4'd2, 5'd0, 1'd1} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd2, 5'd1, 1'd1} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd2, 5'd2, 1'd1} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd2, 5'd3, 1'd1} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd2, 5'd4, 1'd1} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd2, 5'd5, 1'd1} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd2, 5'd6, 1'd1} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd2, 5'd7, 1'd1} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd3, 5'd0, 1'd1} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd3, 5'd1, 1'd1} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd3, 5'd2, 1'd1} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd3, 5'd3, 1'd1} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd3, 5'd4, 1'd1} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd3, 5'd5, 1'd1} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd3, 5'd6, 1'd1} : intpi_lcpll_expected = 4'b0011;
  {PCIE, 4'd3, 5'd7, 1'd1} : intpi_lcpll_expected = 4'b0011;
default: intpi_lcpll_expected = 4'bzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel} )
  {USB, 4'd1, 5'd0, 1'd0} : tx_intpr_expected = 2'b10;
  {USB, 4'd1, 5'd1, 1'd0} : tx_intpr_expected = 2'b10;
  {USB, 4'd1, 5'd2, 1'd0} : tx_intpr_expected = 2'b10;
  {USB, 4'd1, 5'd3, 1'd0} : tx_intpr_expected = 2'b10;
  {USB, 4'd1, 5'd4, 1'd0} : tx_intpr_expected = 2'b10;
  {USB, 4'd1, 5'd5, 1'd0} : tx_intpr_expected = 2'b10;
  {USB, 4'd1, 5'd6, 1'd0} : tx_intpr_expected = 2'b10;
  {USB, 4'd1, 5'd7, 1'd0} : tx_intpr_expected = 2'b10;
  {USB, 4'd2, 5'd0, 1'd0} : tx_intpr_expected = 2'b10;
  {USB, 4'd2, 5'd1, 1'd0} : tx_intpr_expected = 2'b10;
  {USB, 4'd2, 5'd2, 1'd0} : tx_intpr_expected = 2'b10;
  {USB, 4'd2, 5'd3, 1'd0} : tx_intpr_expected = 2'b10;
  {USB, 4'd2, 5'd4, 1'd0} : tx_intpr_expected = 2'b10;
  {USB, 4'd2, 5'd5, 1'd0} : tx_intpr_expected = 2'b10;
  {USB, 4'd2, 5'd6, 1'd0} : tx_intpr_expected = 2'b10;
  {USB, 4'd2, 5'd7, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd0, 5'd0, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd0, 5'd1, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd0, 5'd2, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd0, 5'd3, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd0, 5'd4, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd0, 5'd5, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd0, 5'd6, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd0, 5'd7, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd1, 5'd0, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd1, 5'd1, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd1, 5'd2, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd1, 5'd3, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd1, 5'd4, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd1, 5'd5, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd1, 5'd6, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd1, 5'd7, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd2, 5'd0, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd2, 5'd1, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd2, 5'd2, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd2, 5'd3, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd2, 5'd4, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd2, 5'd5, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd2, 5'd6, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd2, 5'd7, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd3, 5'd0, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd3, 5'd1, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd3, 5'd2, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd3, 5'd3, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd3, 5'd4, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd3, 5'd5, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd3, 5'd6, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd3, 5'd7, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd4, 5'd0, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd4, 5'd1, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd4, 5'd2, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd4, 5'd3, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd4, 5'd4, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd4, 5'd5, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd4, 5'd6, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd4, 5'd7, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd5, 5'd0, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd5, 5'd1, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd5, 5'd2, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd5, 5'd3, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd5, 5'd4, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd5, 5'd5, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd5, 5'd6, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd5, 5'd7, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd6, 5'd0, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd6, 5'd1, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd6, 5'd2, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd6, 5'd3, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd6, 5'd4, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd6, 5'd5, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd6, 5'd6, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd6, 5'd7, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd7, 5'd0, 1'd0} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd7, 5'd1, 1'd0} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd7, 5'd2, 1'd0} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd7, 5'd3, 1'd0} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd7, 5'd4, 1'd0} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd7, 5'd5, 1'd0} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd7, 5'd6, 1'd0} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd7, 5'd7, 1'd0} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd8, 5'd0, 1'd0} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd8, 5'd1, 1'd0} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd8, 5'd2, 1'd0} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd8, 5'd3, 1'd0} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd8, 5'd4, 1'd0} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd8, 5'd5, 1'd0} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd8, 5'd6, 1'd0} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd8, 5'd7, 1'd0} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd9, 5'd0, 1'd0} : tx_intpr_expected = 2'b00;
  {SERDES, 4'd9, 5'd1, 1'd0} : tx_intpr_expected = 2'b00;
  {SERDES, 4'd9, 5'd2, 1'd0} : tx_intpr_expected = 2'b00;
  {SERDES, 4'd9, 5'd3, 1'd0} : tx_intpr_expected = 2'b00;
  {SERDES, 4'd9, 5'd4, 1'd0} : tx_intpr_expected = 2'b00;
  {SERDES, 4'd9, 5'd5, 1'd0} : tx_intpr_expected = 2'b00;
  {SERDES, 4'd9, 5'd6, 1'd0} : tx_intpr_expected = 2'b00;
  {SERDES, 4'd9, 5'd7, 1'd0} : tx_intpr_expected = 2'b00;
  {SERDES, 4'd12, 5'd0, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd12, 5'd1, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd12, 5'd2, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd12, 5'd3, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd12, 5'd4, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd12, 5'd5, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd12, 5'd6, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd12, 5'd7, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd13, 5'd0, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd13, 5'd1, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd13, 5'd2, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd13, 5'd3, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd13, 5'd4, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd13, 5'd5, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd13, 5'd6, 1'd0} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd13, 5'd7, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd0, 5'd0, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd0, 5'd1, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd0, 5'd2, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd0, 5'd3, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd0, 5'd4, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd0, 5'd5, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd0, 5'd6, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd0, 5'd7, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd1, 5'd0, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd1, 5'd1, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd1, 5'd2, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd1, 5'd3, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd1, 5'd4, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd1, 5'd5, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd1, 5'd6, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd1, 5'd7, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd2, 5'd0, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd2, 5'd1, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd2, 5'd2, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd2, 5'd3, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd2, 5'd4, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd2, 5'd5, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd2, 5'd6, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd2, 5'd7, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd3, 5'd0, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd3, 5'd1, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd3, 5'd2, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd3, 5'd3, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd3, 5'd4, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd3, 5'd5, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd3, 5'd6, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd3, 5'd7, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd4, 5'd0, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd4, 5'd1, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd4, 5'd2, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd4, 5'd3, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd4, 5'd4, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd4, 5'd5, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd4, 5'd6, 1'd0} : tx_intpr_expected = 2'b10;
  {SAS, 4'd4, 5'd7, 1'd0} : tx_intpr_expected = 2'b10;
  {PCIE, 4'd2, 5'd0, 1'd0} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd2, 5'd1, 1'd0} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd2, 5'd2, 1'd0} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd2, 5'd3, 1'd0} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd2, 5'd4, 1'd0} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd2, 5'd5, 1'd0} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd2, 5'd6, 1'd0} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd2, 5'd7, 1'd0} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd3, 5'd0, 1'd0} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd3, 5'd1, 1'd0} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd3, 5'd2, 1'd0} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd3, 5'd3, 1'd0} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd3, 5'd4, 1'd0} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd3, 5'd5, 1'd0} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd3, 5'd6, 1'd0} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd3, 5'd7, 1'd0} : tx_intpr_expected = 2'b11;
  {USB, 4'd1, 5'd0, 1'd1} : tx_intpr_expected = 2'b10;
  {USB, 4'd1, 5'd1, 1'd1} : tx_intpr_expected = 2'b10;
  {USB, 4'd1, 5'd2, 1'd1} : tx_intpr_expected = 2'b10;
  {USB, 4'd1, 5'd3, 1'd1} : tx_intpr_expected = 2'b10;
  {USB, 4'd1, 5'd4, 1'd1} : tx_intpr_expected = 2'b10;
  {USB, 4'd1, 5'd5, 1'd1} : tx_intpr_expected = 2'b10;
  {USB, 4'd1, 5'd6, 1'd1} : tx_intpr_expected = 2'b10;
  {USB, 4'd1, 5'd7, 1'd1} : tx_intpr_expected = 2'b10;
  {USB, 4'd2, 5'd0, 1'd1} : tx_intpr_expected = 2'b10;
  {USB, 4'd2, 5'd1, 1'd1} : tx_intpr_expected = 2'b10;
  {USB, 4'd2, 5'd2, 1'd1} : tx_intpr_expected = 2'b10;
  {USB, 4'd2, 5'd3, 1'd1} : tx_intpr_expected = 2'b10;
  {USB, 4'd2, 5'd4, 1'd1} : tx_intpr_expected = 2'b10;
  {USB, 4'd2, 5'd5, 1'd1} : tx_intpr_expected = 2'b10;
  {USB, 4'd2, 5'd6, 1'd1} : tx_intpr_expected = 2'b10;
  {USB, 4'd2, 5'd7, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd0, 5'd0, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd0, 5'd1, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd0, 5'd2, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd0, 5'd3, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd0, 5'd4, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd0, 5'd5, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd0, 5'd6, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd0, 5'd7, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd1, 5'd0, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd1, 5'd1, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd1, 5'd2, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd1, 5'd3, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd1, 5'd4, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd1, 5'd5, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd1, 5'd6, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd1, 5'd7, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd2, 5'd0, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd2, 5'd1, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd2, 5'd2, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd2, 5'd3, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd2, 5'd4, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd2, 5'd5, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd2, 5'd6, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd2, 5'd7, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd3, 5'd0, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd3, 5'd1, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd3, 5'd2, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd3, 5'd3, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd3, 5'd4, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd3, 5'd5, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd3, 5'd6, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd3, 5'd7, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd4, 5'd0, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd4, 5'd1, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd4, 5'd2, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd4, 5'd3, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd4, 5'd4, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd4, 5'd5, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd4, 5'd6, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd4, 5'd7, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd5, 5'd0, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd5, 5'd1, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd5, 5'd2, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd5, 5'd3, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd5, 5'd4, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd5, 5'd5, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd5, 5'd6, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd5, 5'd7, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd6, 5'd0, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd6, 5'd1, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd6, 5'd2, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd6, 5'd3, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd6, 5'd4, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd6, 5'd5, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd6, 5'd6, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd6, 5'd7, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd7, 5'd0, 1'd1} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd7, 5'd1, 1'd1} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd7, 5'd2, 1'd1} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd7, 5'd3, 1'd1} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd7, 5'd4, 1'd1} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd7, 5'd5, 1'd1} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd7, 5'd6, 1'd1} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd7, 5'd7, 1'd1} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd8, 5'd0, 1'd1} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd8, 5'd1, 1'd1} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd8, 5'd2, 1'd1} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd8, 5'd3, 1'd1} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd8, 5'd4, 1'd1} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd8, 5'd5, 1'd1} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd8, 5'd6, 1'd1} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd8, 5'd7, 1'd1} : tx_intpr_expected = 2'b01;
  {SERDES, 4'd9, 5'd0, 1'd1} : tx_intpr_expected = 2'b00;
  {SERDES, 4'd9, 5'd1, 1'd1} : tx_intpr_expected = 2'b00;
  {SERDES, 4'd9, 5'd2, 1'd1} : tx_intpr_expected = 2'b00;
  {SERDES, 4'd9, 5'd3, 1'd1} : tx_intpr_expected = 2'b00;
  {SERDES, 4'd9, 5'd4, 1'd1} : tx_intpr_expected = 2'b00;
  {SERDES, 4'd9, 5'd5, 1'd1} : tx_intpr_expected = 2'b00;
  {SERDES, 4'd9, 5'd6, 1'd1} : tx_intpr_expected = 2'b00;
  {SERDES, 4'd9, 5'd7, 1'd1} : tx_intpr_expected = 2'b00;
  {SERDES, 4'd12, 5'd0, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd12, 5'd1, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd12, 5'd2, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd12, 5'd3, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd12, 5'd4, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd12, 5'd5, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd12, 5'd6, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd12, 5'd7, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd13, 5'd0, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd13, 5'd1, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd13, 5'd2, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd13, 5'd3, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd13, 5'd4, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd13, 5'd5, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd13, 5'd6, 1'd1} : tx_intpr_expected = 2'b10;
  {SERDES, 4'd13, 5'd7, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd0, 5'd0, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd0, 5'd1, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd0, 5'd2, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd0, 5'd3, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd0, 5'd4, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd0, 5'd5, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd0, 5'd6, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd0, 5'd7, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd1, 5'd0, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd1, 5'd1, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd1, 5'd2, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd1, 5'd3, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd1, 5'd4, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd1, 5'd5, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd1, 5'd6, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd1, 5'd7, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd2, 5'd0, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd2, 5'd1, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd2, 5'd2, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd2, 5'd3, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd2, 5'd4, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd2, 5'd5, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd2, 5'd6, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd2, 5'd7, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd3, 5'd0, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd3, 5'd1, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd3, 5'd2, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd3, 5'd3, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd3, 5'd4, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd3, 5'd5, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd3, 5'd6, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd3, 5'd7, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd4, 5'd0, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd4, 5'd1, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd4, 5'd2, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd4, 5'd3, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd4, 5'd4, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd4, 5'd5, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd4, 5'd6, 1'd1} : tx_intpr_expected = 2'b10;
  {SAS, 4'd4, 5'd7, 1'd1} : tx_intpr_expected = 2'b10;
  {PCIE, 4'd2, 5'd0, 1'd1} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd2, 5'd1, 1'd1} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd2, 5'd2, 1'd1} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd2, 5'd3, 1'd1} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd2, 5'd4, 1'd1} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd2, 5'd5, 1'd1} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd2, 5'd6, 1'd1} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd2, 5'd7, 1'd1} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd3, 5'd0, 1'd1} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd3, 5'd1, 1'd1} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd3, 5'd2, 1'd1} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd3, 5'd3, 1'd1} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd3, 5'd4, 1'd1} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd3, 5'd5, 1'd1} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd3, 5'd6, 1'd1} : tx_intpr_expected = 2'b11;
  {PCIE, 4'd3, 5'd7, 1'd1} : tx_intpr_expected = 2'b11;
default: tx_intpr_expected = 2'bzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel} )
  {USB, 4'd1, 5'd0, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd1, 5'd1, 1'd0} : init_txfoffs_expected = 10'b1111011111;
  {USB, 4'd1, 5'd2, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd1, 5'd3, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd1, 5'd4, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd1, 5'd5, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd1, 5'd6, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd1, 5'd7, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd2, 5'd0, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd2, 5'd1, 1'd0} : init_txfoffs_expected = 10'b1111011111;
  {USB, 4'd2, 5'd2, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd2, 5'd3, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd2, 5'd4, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd2, 5'd5, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd2, 5'd6, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd2, 5'd7, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd0, 5'd0, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd0, 5'd1, 1'd0} : init_txfoffs_expected = 10'b1111011111;
  {SERDES, 4'd0, 5'd2, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd0, 5'd3, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd0, 5'd4, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd0, 5'd5, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd0, 5'd6, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd0, 5'd7, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd1, 5'd0, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd1, 5'd1, 1'd0} : init_txfoffs_expected = 10'b0000011010;
  {SERDES, 4'd1, 5'd2, 1'd0} : init_txfoffs_expected = 10'b0000110100;
  {SERDES, 4'd1, 5'd3, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd1, 5'd4, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd1, 5'd5, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd1, 5'd6, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd1, 5'd7, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd2, 5'd0, 1'd0} : init_txfoffs_expected = 10'b0000101000;
  {SERDES, 4'd2, 5'd1, 1'd0} : init_txfoffs_expected = 10'b0000011000;
  {SERDES, 4'd2, 5'd2, 1'd0} : init_txfoffs_expected = 10'b0000011000;
  {SERDES, 4'd2, 5'd3, 1'd0} : init_txfoffs_expected = 10'b1111011000;
  {SERDES, 4'd2, 5'd4, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd2, 5'd5, 1'd0} : init_txfoffs_expected = 10'b1111011000;
  {SERDES, 4'd2, 5'd6, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd2, 5'd7, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd3, 5'd0, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd3, 5'd1, 1'd0} : init_txfoffs_expected = 10'b0000011010;
  {SERDES, 4'd3, 5'd2, 1'd0} : init_txfoffs_expected = 10'b0000110100;
  {SERDES, 4'd3, 5'd3, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd3, 5'd4, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd3, 5'd5, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd3, 5'd6, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd3, 5'd7, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd4, 5'd0, 1'd0} : init_txfoffs_expected = 10'b0000101000;
  {SERDES, 4'd4, 5'd1, 1'd0} : init_txfoffs_expected = 10'b0000011000;
  {SERDES, 4'd4, 5'd2, 1'd0} : init_txfoffs_expected = 10'b0000011000;
  {SERDES, 4'd4, 5'd3, 1'd0} : init_txfoffs_expected = 10'b1111011000;
  {SERDES, 4'd4, 5'd4, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd4, 5'd5, 1'd0} : init_txfoffs_expected = 10'b1111011000;
  {SERDES, 4'd4, 5'd6, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd4, 5'd7, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd5, 5'd0, 1'd0} : init_txfoffs_expected = 10'b0000100010;
  {SERDES, 4'd5, 5'd1, 1'd0} : init_txfoffs_expected = 10'b1111101100;
  {SERDES, 4'd5, 5'd2, 1'd0} : init_txfoffs_expected = 10'b0000100010;
  {SERDES, 4'd5, 5'd3, 1'd0} : init_txfoffs_expected = 10'b0000100010;
  {SERDES, 4'd5, 5'd4, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd5, 5'd5, 1'd0} : init_txfoffs_expected = 10'b0000100010;
  {SERDES, 4'd5, 5'd6, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd5, 5'd7, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd6, 5'd0, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd6, 5'd1, 1'd0} : init_txfoffs_expected = 10'b0000011010;
  {SERDES, 4'd6, 5'd2, 1'd0} : init_txfoffs_expected = 10'b0000110100;
  {SERDES, 4'd6, 5'd3, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd6, 5'd4, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd6, 5'd5, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd6, 5'd6, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd6, 5'd7, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd7, 5'd0, 1'd0} : init_txfoffs_expected = 10'b0000011000;
  {SERDES, 4'd7, 5'd1, 1'd0} : init_txfoffs_expected = 10'b0000011000;
  {SERDES, 4'd7, 5'd2, 1'd0} : init_txfoffs_expected = 10'b1111100101;
  {SERDES, 4'd7, 5'd3, 1'd0} : init_txfoffs_expected = 10'b0000011000;
  {SERDES, 4'd7, 5'd4, 1'd0} : init_txfoffs_expected = 10'b1111011000;
  {SERDES, 4'd7, 5'd5, 1'd0} : init_txfoffs_expected = 10'b0000011000;
  {SERDES, 4'd7, 5'd6, 1'd0} : init_txfoffs_expected = 10'b1111011000;
  {SERDES, 4'd7, 5'd7, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd8, 5'd0, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd8, 5'd1, 1'd0} : init_txfoffs_expected = 10'b1111101000;
  {SERDES, 4'd8, 5'd2, 1'd0} : init_txfoffs_expected = 10'b0000011000;
  {SERDES, 4'd8, 5'd3, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd8, 5'd4, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd8, 5'd5, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd8, 5'd6, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd8, 5'd7, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd9, 5'd0, 1'd0} : init_txfoffs_expected = 10'b0000011101;
  {SERDES, 4'd9, 5'd1, 1'd0} : init_txfoffs_expected = 10'b0000010001;
  {SERDES, 4'd9, 5'd2, 1'd0} : init_txfoffs_expected = 10'b0000101001;
  {SERDES, 4'd9, 5'd3, 1'd0} : init_txfoffs_expected = 10'b1111100011;
  {SERDES, 4'd9, 5'd4, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd9, 5'd5, 1'd0} : init_txfoffs_expected = 10'b1111100011;
  {SERDES, 4'd9, 5'd6, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd9, 5'd7, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd12, 5'd0, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd12, 5'd1, 1'd0} : init_txfoffs_expected = 10'b1111011111;
  {SERDES, 4'd12, 5'd2, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd12, 5'd3, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd12, 5'd4, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd12, 5'd5, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd12, 5'd6, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd12, 5'd7, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd13, 5'd0, 1'd0} : init_txfoffs_expected = 10'b0000101000;
  {SERDES, 4'd13, 5'd1, 1'd0} : init_txfoffs_expected = 10'b0000011000;
  {SERDES, 4'd13, 5'd2, 1'd0} : init_txfoffs_expected = 10'b0000011000;
  {SERDES, 4'd13, 5'd3, 1'd0} : init_txfoffs_expected = 10'b1111011000;
  {SERDES, 4'd13, 5'd4, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd13, 5'd5, 1'd0} : init_txfoffs_expected = 10'b1111011000;
  {SERDES, 4'd13, 5'd6, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd13, 5'd7, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd0, 5'd0, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd0, 5'd1, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd0, 5'd2, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd0, 5'd3, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd0, 5'd4, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd0, 5'd5, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd0, 5'd6, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd0, 5'd7, 1'd0} : init_txfoffs_expected = 10'b1111101011;
  {SAS, 4'd1, 5'd0, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd1, 5'd1, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd1, 5'd2, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd1, 5'd3, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd1, 5'd4, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd1, 5'd5, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd1, 5'd6, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd1, 5'd7, 1'd0} : init_txfoffs_expected = 10'b1111101011;
  {SAS, 4'd2, 5'd0, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd2, 5'd1, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd2, 5'd2, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd2, 5'd3, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd2, 5'd4, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd2, 5'd5, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd2, 5'd6, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd2, 5'd7, 1'd0} : init_txfoffs_expected = 10'b1111101011;
  {SAS, 4'd3, 5'd0, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd3, 5'd1, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd3, 5'd2, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd3, 5'd3, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd3, 5'd4, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd3, 5'd5, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd3, 5'd6, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd3, 5'd7, 1'd0} : init_txfoffs_expected = 10'b1111101011;
  {SAS, 4'd4, 5'd0, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd4, 5'd1, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd4, 5'd2, 1'd0} : init_txfoffs_expected = 10'b1111100011;
  {SAS, 4'd4, 5'd3, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd4, 5'd4, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd4, 5'd5, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd4, 5'd6, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd4, 5'd7, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd2, 5'd0, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd2, 5'd1, 1'd0} : init_txfoffs_expected = 10'b0000101001;
  {PCIE, 4'd2, 5'd2, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd2, 5'd3, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd2, 5'd4, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd2, 5'd5, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd2, 5'd6, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd2, 5'd7, 1'd0} : init_txfoffs_expected = 10'b0000100000;
  {PCIE, 4'd3, 5'd0, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd3, 5'd1, 1'd0} : init_txfoffs_expected = 10'b0000101001;
  {PCIE, 4'd3, 5'd2, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd3, 5'd3, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd3, 5'd4, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd3, 5'd5, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd3, 5'd6, 1'd0} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd3, 5'd7, 1'd0} : init_txfoffs_expected = 10'b0000100000;
  {USB, 4'd1, 5'd0, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd1, 5'd1, 1'd1} : init_txfoffs_expected = 10'b1101111101;
  {USB, 4'd1, 5'd2, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd1, 5'd3, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd1, 5'd4, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd1, 5'd5, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd1, 5'd6, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd1, 5'd7, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd2, 5'd0, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd2, 5'd1, 1'd1} : init_txfoffs_expected = 10'b1101111101;
  {USB, 4'd2, 5'd2, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd2, 5'd3, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd2, 5'd4, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd2, 5'd5, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd2, 5'd6, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {USB, 4'd2, 5'd7, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd0, 5'd0, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd0, 5'd1, 1'd1} : init_txfoffs_expected = 10'b1101111101;
  {SERDES, 4'd0, 5'd2, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd0, 5'd3, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd0, 5'd4, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd0, 5'd5, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd0, 5'd6, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd0, 5'd7, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd1, 5'd0, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd1, 5'd1, 1'd1} : init_txfoffs_expected = 10'b1111001100;
  {SERDES, 4'd1, 5'd2, 1'd1} : init_txfoffs_expected = 10'b1111001100;
  {SERDES, 4'd1, 5'd3, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd1, 5'd4, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd1, 5'd5, 1'd1} : init_txfoffs_expected = 10'b0001010111;
  {SERDES, 4'd1, 5'd6, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd1, 5'd7, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd2, 5'd0, 1'd1} : init_txfoffs_expected = 10'b1111011000;
  {SERDES, 4'd2, 5'd1, 1'd1} : init_txfoffs_expected = 10'b0000011000;
  {SERDES, 4'd2, 5'd2, 1'd1} : init_txfoffs_expected = 10'b1111000011;
  {SERDES, 4'd2, 5'd3, 1'd1} : init_txfoffs_expected = 10'b1111011000;
  {SERDES, 4'd2, 5'd4, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd2, 5'd5, 1'd1} : init_txfoffs_expected = 10'b1111011000;
  {SERDES, 4'd2, 5'd6, 1'd1} : init_txfoffs_expected = 10'b0001000010;
  {SERDES, 4'd2, 5'd7, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd3, 5'd0, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd3, 5'd1, 1'd1} : init_txfoffs_expected = 10'b1111001100;
  {SERDES, 4'd3, 5'd2, 1'd1} : init_txfoffs_expected = 10'b1111001100;
  {SERDES, 4'd3, 5'd3, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd3, 5'd4, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd3, 5'd5, 1'd1} : init_txfoffs_expected = 10'b0001010111;
  {SERDES, 4'd3, 5'd6, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd3, 5'd7, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd4, 5'd0, 1'd1} : init_txfoffs_expected = 10'b1111011000;
  {SERDES, 4'd4, 5'd1, 1'd1} : init_txfoffs_expected = 10'b0000011000;
  {SERDES, 4'd4, 5'd2, 1'd1} : init_txfoffs_expected = 10'b1111000011;
  {SERDES, 4'd4, 5'd3, 1'd1} : init_txfoffs_expected = 10'b1111011000;
  {SERDES, 4'd4, 5'd4, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd4, 5'd5, 1'd1} : init_txfoffs_expected = 10'b1111011000;
  {SERDES, 4'd4, 5'd6, 1'd1} : init_txfoffs_expected = 10'b0001000010;
  {SERDES, 4'd4, 5'd7, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd5, 5'd0, 1'd1} : init_txfoffs_expected = 10'b0000100010;
  {SERDES, 4'd5, 5'd1, 1'd1} : init_txfoffs_expected = 10'b1111101100;
  {SERDES, 4'd5, 5'd2, 1'd1} : init_txfoffs_expected = 10'b1110110110;
  {SERDES, 4'd5, 5'd3, 1'd1} : init_txfoffs_expected = 10'b0000100010;
  {SERDES, 4'd5, 5'd4, 1'd1} : init_txfoffs_expected = 10'b0010101000;
  {SERDES, 4'd5, 5'd5, 1'd1} : init_txfoffs_expected = 10'b0000100010;
  {SERDES, 4'd5, 5'd6, 1'd1} : init_txfoffs_expected = 10'b0010101000;
  {SERDES, 4'd5, 5'd7, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd6, 5'd0, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd6, 5'd1, 1'd1} : init_txfoffs_expected = 10'b1111001100;
  {SERDES, 4'd6, 5'd2, 1'd1} : init_txfoffs_expected = 10'b1111001100;
  {SERDES, 4'd6, 5'd3, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd6, 5'd4, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd6, 5'd5, 1'd1} : init_txfoffs_expected = 10'b0001010111;
  {SERDES, 4'd6, 5'd6, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd6, 5'd7, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd7, 5'd0, 1'd1} : init_txfoffs_expected = 10'b0000011000;
  {SERDES, 4'd7, 5'd1, 1'd1} : init_txfoffs_expected = 10'b1101111111;
  {SERDES, 4'd7, 5'd2, 1'd1} : init_txfoffs_expected = 10'b0010110000;
  {SERDES, 4'd7, 5'd3, 1'd1} : init_txfoffs_expected = 10'b0000011000;
  {SERDES, 4'd7, 5'd4, 1'd1} : init_txfoffs_expected = 10'b0001000010;
  {SERDES, 4'd7, 5'd5, 1'd1} : init_txfoffs_expected = 10'b0001101101;
  {SERDES, 4'd7, 5'd6, 1'd1} : init_txfoffs_expected = 10'b0000011000;
  {SERDES, 4'd7, 5'd7, 1'd1} : init_txfoffs_expected = 10'b0001000010;
  {SERDES, 4'd8, 5'd0, 1'd1} : init_txfoffs_expected = 10'b0001110111;
  {SERDES, 4'd8, 5'd1, 1'd1} : init_txfoffs_expected = 10'b1111101000;
  {SERDES, 4'd8, 5'd2, 1'd1} : init_txfoffs_expected = 10'b0000011000;
  {SERDES, 4'd8, 5'd3, 1'd1} : init_txfoffs_expected = 10'b0001110111;
  {SERDES, 4'd8, 5'd4, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd8, 5'd5, 1'd1} : init_txfoffs_expected = 10'b0001110111;
  {SERDES, 4'd8, 5'd6, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd8, 5'd7, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd9, 5'd0, 1'd1} : init_txfoffs_expected = 10'b0001010111;
  {SERDES, 4'd9, 5'd1, 1'd1} : init_txfoffs_expected = 10'b1111001100;
  {SERDES, 4'd9, 5'd2, 1'd1} : init_txfoffs_expected = 10'b0000101001;
  {SERDES, 4'd9, 5'd3, 1'd1} : init_txfoffs_expected = 10'b1101101110;
  {SERDES, 4'd9, 5'd4, 1'd1} : init_txfoffs_expected = 10'b1101101110;
  {SERDES, 4'd9, 5'd5, 1'd1} : init_txfoffs_expected = 10'b1101101110;
  {SERDES, 4'd9, 5'd6, 1'd1} : init_txfoffs_expected = 10'b1101101110;
  {SERDES, 4'd9, 5'd7, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd12, 5'd0, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd12, 5'd1, 1'd1} : init_txfoffs_expected = 10'b1101111101;
  {SERDES, 4'd12, 5'd2, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd12, 5'd3, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd12, 5'd4, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd12, 5'd5, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd12, 5'd6, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd12, 5'd7, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd13, 5'd0, 1'd1} : init_txfoffs_expected = 10'b1111011000;
  {SERDES, 4'd13, 5'd1, 1'd1} : init_txfoffs_expected = 10'b0000011000;
  {SERDES, 4'd13, 5'd2, 1'd1} : init_txfoffs_expected = 10'b1111000011;
  {SERDES, 4'd13, 5'd3, 1'd1} : init_txfoffs_expected = 10'b1111011000;
  {SERDES, 4'd13, 5'd4, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SERDES, 4'd13, 5'd5, 1'd1} : init_txfoffs_expected = 10'b1111011000;
  {SERDES, 4'd13, 5'd6, 1'd1} : init_txfoffs_expected = 10'b0001000010;
  {SERDES, 4'd13, 5'd7, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd0, 5'd0, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd0, 5'd1, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd0, 5'd2, 1'd1} : init_txfoffs_expected = 10'b0010010010;
  {SAS, 4'd0, 5'd3, 1'd1} : init_txfoffs_expected = 10'b0010110101;
  {SAS, 4'd0, 5'd4, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd0, 5'd5, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd0, 5'd6, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd0, 5'd7, 1'd1} : init_txfoffs_expected = 10'b0001010101;
  {SAS, 4'd1, 5'd0, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd1, 5'd1, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd1, 5'd2, 1'd1} : init_txfoffs_expected = 10'b0010010010;
  {SAS, 4'd1, 5'd3, 1'd1} : init_txfoffs_expected = 10'b0010110101;
  {SAS, 4'd1, 5'd4, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd1, 5'd5, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd1, 5'd6, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd1, 5'd7, 1'd1} : init_txfoffs_expected = 10'b0001010101;
  {SAS, 4'd2, 5'd0, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd2, 5'd1, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd2, 5'd2, 1'd1} : init_txfoffs_expected = 10'b0010010010;
  {SAS, 4'd2, 5'd3, 1'd1} : init_txfoffs_expected = 10'b0010110101;
  {SAS, 4'd2, 5'd4, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd2, 5'd5, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd2, 5'd6, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd2, 5'd7, 1'd1} : init_txfoffs_expected = 10'b0001010101;
  {SAS, 4'd3, 5'd0, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd3, 5'd1, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd3, 5'd2, 1'd1} : init_txfoffs_expected = 10'b0010010010;
  {SAS, 4'd3, 5'd3, 1'd1} : init_txfoffs_expected = 10'b0010110101;
  {SAS, 4'd3, 5'd4, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd3, 5'd5, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd3, 5'd6, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd3, 5'd7, 1'd1} : init_txfoffs_expected = 10'b0001010101;
  {SAS, 4'd4, 5'd0, 1'd1} : init_txfoffs_expected = 10'b0010010010;
  {SAS, 4'd4, 5'd1, 1'd1} : init_txfoffs_expected = 10'b0001010111;
  {SAS, 4'd4, 5'd2, 1'd1} : init_txfoffs_expected = 10'b1101101110;
  {SAS, 4'd4, 5'd3, 1'd1} : init_txfoffs_expected = 10'b1101101110;
  {SAS, 4'd4, 5'd4, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd4, 5'd5, 1'd1} : init_txfoffs_expected = 10'b1101101110;
  {SAS, 4'd4, 5'd6, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {SAS, 4'd4, 5'd7, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd2, 5'd0, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd2, 5'd1, 1'd1} : init_txfoffs_expected = 10'b1110101110;
  {PCIE, 4'd2, 5'd2, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd2, 5'd3, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd2, 5'd4, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd2, 5'd5, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd2, 5'd6, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd2, 5'd7, 1'd1} : init_txfoffs_expected = 10'b1110000000;
  {PCIE, 4'd3, 5'd0, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd3, 5'd1, 1'd1} : init_txfoffs_expected = 10'b1110101110;
  {PCIE, 4'd3, 5'd2, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd3, 5'd3, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd3, 5'd4, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd3, 5'd5, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd3, 5'd6, 1'd1} : init_txfoffs_expected = 10'b0000000000;
  {PCIE, 4'd3, 5'd7, 1'd1} : init_txfoffs_expected = 10'b1110000000;
default: init_txfoffs_expected = 10'bzzzzzzzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel} )
  {USB, 4'd1, 5'd0, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd1, 5'd1, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd1, 5'd2, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd1, 5'd3, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd1, 5'd4, 1'd0} : speed_thresh_expected = 12'b011111100000;
  {USB, 4'd1, 5'd5, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd1, 5'd6, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd1, 5'd7, 1'd0} : speed_thresh_expected = 12'b011111011010;
  {USB, 4'd2, 5'd0, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd2, 5'd1, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd2, 5'd2, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd2, 5'd3, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd2, 5'd4, 1'd0} : speed_thresh_expected = 12'b011111100000;
  {USB, 4'd2, 5'd5, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd2, 5'd6, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd2, 5'd7, 1'd0} : speed_thresh_expected = 12'b011111011010;
  {SERDES, 4'd0, 5'd0, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd0, 5'd1, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd0, 5'd2, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd0, 5'd3, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd0, 5'd4, 1'd0} : speed_thresh_expected = 12'b011111100000;
  {SERDES, 4'd0, 5'd5, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd0, 5'd6, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd0, 5'd7, 1'd0} : speed_thresh_expected = 12'b011111011010;
  {SERDES, 4'd1, 5'd0, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd1, 5'd1, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd1, 5'd2, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd1, 5'd3, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd1, 5'd4, 1'd0} : speed_thresh_expected = 12'b011111100000;
  {SERDES, 4'd1, 5'd5, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd1, 5'd6, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd1, 5'd7, 1'd0} : speed_thresh_expected = 12'b011111011010;
  {SERDES, 4'd2, 5'd0, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd2, 5'd1, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd2, 5'd2, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd2, 5'd3, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd2, 5'd4, 1'd0} : speed_thresh_expected = 12'b011110111100;
  {SERDES, 4'd2, 5'd5, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd2, 5'd6, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd2, 5'd7, 1'd0} : speed_thresh_expected = 12'b011110110110;
  {SERDES, 4'd3, 5'd0, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd3, 5'd1, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd3, 5'd2, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd3, 5'd3, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd3, 5'd4, 1'd0} : speed_thresh_expected = 12'b011111100000;
  {SERDES, 4'd3, 5'd5, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd3, 5'd6, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd3, 5'd7, 1'd0} : speed_thresh_expected = 12'b011111011010;
  {SERDES, 4'd4, 5'd0, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd4, 5'd1, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd4, 5'd2, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd4, 5'd3, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd4, 5'd4, 1'd0} : speed_thresh_expected = 12'b011110111100;
  {SERDES, 4'd4, 5'd5, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd4, 5'd6, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd4, 5'd7, 1'd0} : speed_thresh_expected = 12'b011110110110;
  {SERDES, 4'd5, 5'd0, 1'd0} : speed_thresh_expected = 12'b011111101111;
  {SERDES, 4'd5, 5'd1, 1'd0} : speed_thresh_expected = 12'b011111101111;
  {SERDES, 4'd5, 5'd2, 1'd0} : speed_thresh_expected = 12'b011111101111;
  {SERDES, 4'd5, 5'd3, 1'd0} : speed_thresh_expected = 12'b011111101111;
  {SERDES, 4'd5, 5'd4, 1'd0} : speed_thresh_expected = 12'b100000000000;
  {SERDES, 4'd5, 5'd5, 1'd0} : speed_thresh_expected = 12'b011111101111;
  {SERDES, 4'd5, 5'd6, 1'd0} : speed_thresh_expected = 12'b011111101111;
  {SERDES, 4'd5, 5'd7, 1'd0} : speed_thresh_expected = 12'b011111111001;
  {SERDES, 4'd6, 5'd0, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd6, 5'd1, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd6, 5'd2, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd6, 5'd3, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd6, 5'd4, 1'd0} : speed_thresh_expected = 12'b011111100000;
  {SERDES, 4'd6, 5'd5, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd6, 5'd6, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd6, 5'd7, 1'd0} : speed_thresh_expected = 12'b011111011010;
  {SERDES, 4'd7, 5'd0, 1'd0} : speed_thresh_expected = 12'b011110111111;
  {SERDES, 4'd7, 5'd1, 1'd0} : speed_thresh_expected = 12'b011110111111;
  {SERDES, 4'd7, 5'd2, 1'd0} : speed_thresh_expected = 12'b011110111111;
  {SERDES, 4'd7, 5'd3, 1'd0} : speed_thresh_expected = 12'b011110111111;
  {SERDES, 4'd7, 5'd4, 1'd0} : speed_thresh_expected = 12'b011111001111;
  {SERDES, 4'd7, 5'd5, 1'd0} : speed_thresh_expected = 12'b011110111111;
  {SERDES, 4'd7, 5'd6, 1'd0} : speed_thresh_expected = 12'b011110111111;
  {SERDES, 4'd7, 5'd7, 1'd0} : speed_thresh_expected = 12'b011111001001;
  {SERDES, 4'd8, 5'd0, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd8, 5'd1, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd8, 5'd2, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd8, 5'd3, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd8, 5'd4, 1'd0} : speed_thresh_expected = 12'b011110111100;
  {SERDES, 4'd8, 5'd5, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd8, 5'd6, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd8, 5'd7, 1'd0} : speed_thresh_expected = 12'b011110110110;
  {SERDES, 4'd9, 5'd0, 1'd0} : speed_thresh_expected = 12'b011111011001;
  {SERDES, 4'd9, 5'd1, 1'd0} : speed_thresh_expected = 12'b011111011001;
  {SERDES, 4'd9, 5'd2, 1'd0} : speed_thresh_expected = 12'b011111011001;
  {SERDES, 4'd9, 5'd3, 1'd0} : speed_thresh_expected = 12'b011111011001;
  {SERDES, 4'd9, 5'd4, 1'd0} : speed_thresh_expected = 12'b011111101001;
  {SERDES, 4'd9, 5'd5, 1'd0} : speed_thresh_expected = 12'b011111011001;
  {SERDES, 4'd9, 5'd6, 1'd0} : speed_thresh_expected = 12'b011111011001;
  {SERDES, 4'd9, 5'd7, 1'd0} : speed_thresh_expected = 12'b011111100011;
  {SERDES, 4'd12, 5'd0, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd12, 5'd1, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd12, 5'd2, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd12, 5'd3, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd12, 5'd4, 1'd0} : speed_thresh_expected = 12'b011111100000;
  {SERDES, 4'd12, 5'd5, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd12, 5'd6, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd12, 5'd7, 1'd0} : speed_thresh_expected = 12'b011111011010;
  {SERDES, 4'd13, 5'd0, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd13, 5'd1, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd13, 5'd2, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd13, 5'd3, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd13, 5'd4, 1'd0} : speed_thresh_expected = 12'b011110111100;
  {SERDES, 4'd13, 5'd5, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd13, 5'd6, 1'd0} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd13, 5'd7, 1'd0} : speed_thresh_expected = 12'b011110110110;
  {SAS, 4'd0, 5'd0, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd0, 5'd1, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd0, 5'd2, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd0, 5'd3, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd0, 5'd4, 1'd0} : speed_thresh_expected = 12'b011111100000;
  {SAS, 4'd0, 5'd5, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd0, 5'd6, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd0, 5'd7, 1'd0} : speed_thresh_expected = 12'b011111011010;
  {SAS, 4'd1, 5'd0, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd1, 5'd1, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd1, 5'd2, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd1, 5'd3, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd1, 5'd4, 1'd0} : speed_thresh_expected = 12'b011111100000;
  {SAS, 4'd1, 5'd5, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd1, 5'd6, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd1, 5'd7, 1'd0} : speed_thresh_expected = 12'b011111011010;
  {SAS, 4'd2, 5'd0, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd2, 5'd1, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd2, 5'd2, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd2, 5'd3, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd2, 5'd4, 1'd0} : speed_thresh_expected = 12'b011111100000;
  {SAS, 4'd2, 5'd5, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd2, 5'd6, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd2, 5'd7, 1'd0} : speed_thresh_expected = 12'b011111011010;
  {SAS, 4'd3, 5'd0, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd3, 5'd1, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd3, 5'd2, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd3, 5'd3, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd3, 5'd4, 1'd0} : speed_thresh_expected = 12'b011111100000;
  {SAS, 4'd3, 5'd5, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd3, 5'd6, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd3, 5'd7, 1'd0} : speed_thresh_expected = 12'b011111011010;
  {SAS, 4'd4, 5'd0, 1'd0} : speed_thresh_expected = 12'b011110100101;
  {SAS, 4'd4, 5'd1, 1'd0} : speed_thresh_expected = 12'b011110100101;
  {SAS, 4'd4, 5'd2, 1'd0} : speed_thresh_expected = 12'b011110100101;
  {SAS, 4'd4, 5'd3, 1'd0} : speed_thresh_expected = 12'b011110100101;
  {SAS, 4'd4, 5'd4, 1'd0} : speed_thresh_expected = 12'b011110110100;
  {SAS, 4'd4, 5'd5, 1'd0} : speed_thresh_expected = 12'b011110100101;
  {SAS, 4'd4, 5'd6, 1'd0} : speed_thresh_expected = 12'b011110100101;
  {SAS, 4'd4, 5'd7, 1'd0} : speed_thresh_expected = 12'b011110101110;
  {PCIE, 4'd2, 5'd0, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd2, 5'd1, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd2, 5'd2, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd2, 5'd3, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd2, 5'd4, 1'd0} : speed_thresh_expected = 12'b011111100000;
  {PCIE, 4'd2, 5'd5, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd2, 5'd6, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd2, 5'd7, 1'd0} : speed_thresh_expected = 12'b011111011010;
  {PCIE, 4'd3, 5'd0, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd3, 5'd1, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd3, 5'd2, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd3, 5'd3, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd3, 5'd4, 1'd0} : speed_thresh_expected = 12'b011111100000;
  {PCIE, 4'd3, 5'd5, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd3, 5'd6, 1'd0} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd3, 5'd7, 1'd0} : speed_thresh_expected = 12'b011111011010;
  {USB, 4'd1, 5'd0, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd1, 5'd1, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd1, 5'd2, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd1, 5'd3, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd1, 5'd4, 1'd1} : speed_thresh_expected = 12'b011111100000;
  {USB, 4'd1, 5'd5, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd1, 5'd6, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd1, 5'd7, 1'd1} : speed_thresh_expected = 12'b011111011010;
  {USB, 4'd2, 5'd0, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd2, 5'd1, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd2, 5'd2, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd2, 5'd3, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd2, 5'd4, 1'd1} : speed_thresh_expected = 12'b011111100000;
  {USB, 4'd2, 5'd5, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd2, 5'd6, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {USB, 4'd2, 5'd7, 1'd1} : speed_thresh_expected = 12'b011111011010;
  {SERDES, 4'd0, 5'd0, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd0, 5'd1, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd0, 5'd2, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd0, 5'd3, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd0, 5'd4, 1'd1} : speed_thresh_expected = 12'b011111100000;
  {SERDES, 4'd0, 5'd5, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd0, 5'd6, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd0, 5'd7, 1'd1} : speed_thresh_expected = 12'b011111011010;
  {SERDES, 4'd1, 5'd0, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd1, 5'd1, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd1, 5'd2, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd1, 5'd3, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd1, 5'd4, 1'd1} : speed_thresh_expected = 12'b011111100000;
  {SERDES, 4'd1, 5'd5, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd1, 5'd6, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd1, 5'd7, 1'd1} : speed_thresh_expected = 12'b011111011010;
  {SERDES, 4'd2, 5'd0, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd2, 5'd1, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd2, 5'd2, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd2, 5'd3, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd2, 5'd4, 1'd1} : speed_thresh_expected = 12'b011110111100;
  {SERDES, 4'd2, 5'd5, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd2, 5'd6, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd2, 5'd7, 1'd1} : speed_thresh_expected = 12'b011110110110;
  {SERDES, 4'd3, 5'd0, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd3, 5'd1, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd3, 5'd2, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd3, 5'd3, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd3, 5'd4, 1'd1} : speed_thresh_expected = 12'b011111100000;
  {SERDES, 4'd3, 5'd5, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd3, 5'd6, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd3, 5'd7, 1'd1} : speed_thresh_expected = 12'b011111011010;
  {SERDES, 4'd4, 5'd0, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd4, 5'd1, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd4, 5'd2, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd4, 5'd3, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd4, 5'd4, 1'd1} : speed_thresh_expected = 12'b011110111100;
  {SERDES, 4'd4, 5'd5, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd4, 5'd6, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd4, 5'd7, 1'd1} : speed_thresh_expected = 12'b011110110110;
  {SERDES, 4'd5, 5'd0, 1'd1} : speed_thresh_expected = 12'b011111101111;
  {SERDES, 4'd5, 5'd1, 1'd1} : speed_thresh_expected = 12'b011111101111;
  {SERDES, 4'd5, 5'd2, 1'd1} : speed_thresh_expected = 12'b011111101111;
  {SERDES, 4'd5, 5'd3, 1'd1} : speed_thresh_expected = 12'b011111101111;
  {SERDES, 4'd5, 5'd4, 1'd1} : speed_thresh_expected = 12'b100000000000;
  {SERDES, 4'd5, 5'd5, 1'd1} : speed_thresh_expected = 12'b011111101111;
  {SERDES, 4'd5, 5'd6, 1'd1} : speed_thresh_expected = 12'b011111101111;
  {SERDES, 4'd5, 5'd7, 1'd1} : speed_thresh_expected = 12'b011111111001;
  {SERDES, 4'd6, 5'd0, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd6, 5'd1, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd6, 5'd2, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd6, 5'd3, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd6, 5'd4, 1'd1} : speed_thresh_expected = 12'b011111100000;
  {SERDES, 4'd6, 5'd5, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd6, 5'd6, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd6, 5'd7, 1'd1} : speed_thresh_expected = 12'b011111011010;
  {SERDES, 4'd7, 5'd0, 1'd1} : speed_thresh_expected = 12'b011110111111;
  {SERDES, 4'd7, 5'd1, 1'd1} : speed_thresh_expected = 12'b011110111111;
  {SERDES, 4'd7, 5'd2, 1'd1} : speed_thresh_expected = 12'b011110111111;
  {SERDES, 4'd7, 5'd3, 1'd1} : speed_thresh_expected = 12'b011110111111;
  {SERDES, 4'd7, 5'd4, 1'd1} : speed_thresh_expected = 12'b011111001111;
  {SERDES, 4'd7, 5'd5, 1'd1} : speed_thresh_expected = 12'b011110111111;
  {SERDES, 4'd7, 5'd6, 1'd1} : speed_thresh_expected = 12'b011110111111;
  {SERDES, 4'd7, 5'd7, 1'd1} : speed_thresh_expected = 12'b011111001001;
  {SERDES, 4'd8, 5'd0, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd8, 5'd1, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd8, 5'd2, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd8, 5'd3, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd8, 5'd4, 1'd1} : speed_thresh_expected = 12'b011110111100;
  {SERDES, 4'd8, 5'd5, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd8, 5'd6, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd8, 5'd7, 1'd1} : speed_thresh_expected = 12'b011110110110;
  {SERDES, 4'd9, 5'd0, 1'd1} : speed_thresh_expected = 12'b011111011001;
  {SERDES, 4'd9, 5'd1, 1'd1} : speed_thresh_expected = 12'b011111011001;
  {SERDES, 4'd9, 5'd2, 1'd1} : speed_thresh_expected = 12'b011111011001;
  {SERDES, 4'd9, 5'd3, 1'd1} : speed_thresh_expected = 12'b011111011001;
  {SERDES, 4'd9, 5'd4, 1'd1} : speed_thresh_expected = 12'b011111101001;
  {SERDES, 4'd9, 5'd5, 1'd1} : speed_thresh_expected = 12'b011111011001;
  {SERDES, 4'd9, 5'd6, 1'd1} : speed_thresh_expected = 12'b011111011001;
  {SERDES, 4'd9, 5'd7, 1'd1} : speed_thresh_expected = 12'b011111100011;
  {SERDES, 4'd12, 5'd0, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd12, 5'd1, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd12, 5'd2, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd12, 5'd3, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd12, 5'd4, 1'd1} : speed_thresh_expected = 12'b011111100000;
  {SERDES, 4'd12, 5'd5, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd12, 5'd6, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SERDES, 4'd12, 5'd7, 1'd1} : speed_thresh_expected = 12'b011111011010;
  {SERDES, 4'd13, 5'd0, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd13, 5'd1, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd13, 5'd2, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd13, 5'd3, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd13, 5'd4, 1'd1} : speed_thresh_expected = 12'b011110111100;
  {SERDES, 4'd13, 5'd5, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd13, 5'd6, 1'd1} : speed_thresh_expected = 12'b011110101100;
  {SERDES, 4'd13, 5'd7, 1'd1} : speed_thresh_expected = 12'b011110110110;
  {SAS, 4'd0, 5'd0, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd0, 5'd1, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd0, 5'd2, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd0, 5'd3, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd0, 5'd4, 1'd1} : speed_thresh_expected = 12'b011111100000;
  {SAS, 4'd0, 5'd5, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd0, 5'd6, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd0, 5'd7, 1'd1} : speed_thresh_expected = 12'b011111011010;
  {SAS, 4'd1, 5'd0, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd1, 5'd1, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd1, 5'd2, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd1, 5'd3, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd1, 5'd4, 1'd1} : speed_thresh_expected = 12'b011111100000;
  {SAS, 4'd1, 5'd5, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd1, 5'd6, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd1, 5'd7, 1'd1} : speed_thresh_expected = 12'b011111011010;
  {SAS, 4'd2, 5'd0, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd2, 5'd1, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd2, 5'd2, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd2, 5'd3, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd2, 5'd4, 1'd1} : speed_thresh_expected = 12'b011111100000;
  {SAS, 4'd2, 5'd5, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd2, 5'd6, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd2, 5'd7, 1'd1} : speed_thresh_expected = 12'b011111011010;
  {SAS, 4'd3, 5'd0, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd3, 5'd1, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd3, 5'd2, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd3, 5'd3, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd3, 5'd4, 1'd1} : speed_thresh_expected = 12'b011111100000;
  {SAS, 4'd3, 5'd5, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd3, 5'd6, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {SAS, 4'd3, 5'd7, 1'd1} : speed_thresh_expected = 12'b011111011010;
  {SAS, 4'd4, 5'd0, 1'd1} : speed_thresh_expected = 12'b011110100101;
  {SAS, 4'd4, 5'd1, 1'd1} : speed_thresh_expected = 12'b011110100101;
  {SAS, 4'd4, 5'd2, 1'd1} : speed_thresh_expected = 12'b011110100101;
  {SAS, 4'd4, 5'd3, 1'd1} : speed_thresh_expected = 12'b011110100101;
  {SAS, 4'd4, 5'd4, 1'd1} : speed_thresh_expected = 12'b011110110100;
  {SAS, 4'd4, 5'd5, 1'd1} : speed_thresh_expected = 12'b011110100101;
  {SAS, 4'd4, 5'd6, 1'd1} : speed_thresh_expected = 12'b011110100101;
  {SAS, 4'd4, 5'd7, 1'd1} : speed_thresh_expected = 12'b011110101110;
  {PCIE, 4'd2, 5'd0, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd2, 5'd1, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd2, 5'd2, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd2, 5'd3, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd2, 5'd4, 1'd1} : speed_thresh_expected = 12'b011111100000;
  {PCIE, 4'd2, 5'd5, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd2, 5'd6, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd2, 5'd7, 1'd1} : speed_thresh_expected = 12'b011111011010;
  {PCIE, 4'd3, 5'd0, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd3, 5'd1, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd3, 5'd2, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd3, 5'd3, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd3, 5'd4, 1'd1} : speed_thresh_expected = 12'b011111100000;
  {PCIE, 4'd3, 5'd5, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd3, 5'd6, 1'd1} : speed_thresh_expected = 12'b011111010000;
  {PCIE, 4'd3, 5'd7, 1'd1} : speed_thresh_expected = 12'b011111011010;
default: speed_thresh_expected = 12'bzzzzzzzzzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel} )
  {USB, 4'd1, 5'd0, 1'd0} : lccap_usb_expected = 1'b0;
  {USB, 4'd1, 5'd1, 1'd0} : lccap_usb_expected = 1'b0;
  {USB, 4'd1, 5'd2, 1'd0} : lccap_usb_expected = 1'b0;
  {USB, 4'd1, 5'd3, 1'd0} : lccap_usb_expected = 1'b0;
  {USB, 4'd1, 5'd4, 1'd0} : lccap_usb_expected = 1'b0;
  {USB, 4'd1, 5'd5, 1'd0} : lccap_usb_expected = 1'b0;
  {USB, 4'd1, 5'd6, 1'd0} : lccap_usb_expected = 1'b0;
  {USB, 4'd1, 5'd7, 1'd0} : lccap_usb_expected = 1'b0;
  {USB, 4'd2, 5'd0, 1'd0} : lccap_usb_expected = 1'b0;
  {USB, 4'd2, 5'd1, 1'd0} : lccap_usb_expected = 1'b0;
  {USB, 4'd2, 5'd2, 1'd0} : lccap_usb_expected = 1'b0;
  {USB, 4'd2, 5'd3, 1'd0} : lccap_usb_expected = 1'b0;
  {USB, 4'd2, 5'd4, 1'd0} : lccap_usb_expected = 1'b0;
  {USB, 4'd2, 5'd5, 1'd0} : lccap_usb_expected = 1'b0;
  {USB, 4'd2, 5'd6, 1'd0} : lccap_usb_expected = 1'b0;
  {USB, 4'd2, 5'd7, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd0, 5'd0, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd0, 5'd1, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd0, 5'd2, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd0, 5'd3, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd0, 5'd4, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd0, 5'd5, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd0, 5'd6, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd0, 5'd7, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd1, 5'd0, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd1, 5'd1, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd1, 5'd2, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd1, 5'd3, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd1, 5'd4, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd1, 5'd5, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd1, 5'd6, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd1, 5'd7, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd2, 5'd0, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd2, 5'd1, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd2, 5'd2, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd2, 5'd3, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd2, 5'd4, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd2, 5'd5, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd2, 5'd6, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd2, 5'd7, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd3, 5'd0, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd3, 5'd1, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd3, 5'd2, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd3, 5'd3, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd3, 5'd4, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd3, 5'd5, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd3, 5'd6, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd3, 5'd7, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd4, 5'd0, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd4, 5'd1, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd4, 5'd2, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd4, 5'd3, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd4, 5'd4, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd4, 5'd5, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd4, 5'd6, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd4, 5'd7, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd5, 5'd0, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd5, 5'd1, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd5, 5'd2, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd5, 5'd3, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd5, 5'd4, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd5, 5'd5, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd5, 5'd6, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd5, 5'd7, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd6, 5'd0, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd6, 5'd1, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd6, 5'd2, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd6, 5'd3, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd6, 5'd4, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd6, 5'd5, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd6, 5'd6, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd6, 5'd7, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd7, 5'd0, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd7, 5'd1, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd7, 5'd2, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd7, 5'd3, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd7, 5'd4, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd7, 5'd5, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd7, 5'd6, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd7, 5'd7, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd8, 5'd0, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd8, 5'd1, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd8, 5'd2, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd8, 5'd3, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd8, 5'd4, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd8, 5'd5, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd8, 5'd6, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd8, 5'd7, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd9, 5'd0, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd9, 5'd1, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd9, 5'd2, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd9, 5'd3, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd9, 5'd4, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd9, 5'd5, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd9, 5'd6, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd9, 5'd7, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd12, 5'd0, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd12, 5'd1, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd12, 5'd2, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd12, 5'd3, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd12, 5'd4, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd12, 5'd5, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd12, 5'd6, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd12, 5'd7, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd13, 5'd0, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd13, 5'd1, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd13, 5'd2, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd13, 5'd3, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd13, 5'd4, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd13, 5'd5, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd13, 5'd6, 1'd0} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd13, 5'd7, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd0, 5'd0, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd0, 5'd1, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd0, 5'd2, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd0, 5'd3, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd0, 5'd4, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd0, 5'd5, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd0, 5'd6, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd0, 5'd7, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd1, 5'd0, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd1, 5'd1, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd1, 5'd2, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd1, 5'd3, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd1, 5'd4, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd1, 5'd5, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd1, 5'd6, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd1, 5'd7, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd2, 5'd0, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd2, 5'd1, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd2, 5'd2, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd2, 5'd3, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd2, 5'd4, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd2, 5'd5, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd2, 5'd6, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd2, 5'd7, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd3, 5'd0, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd3, 5'd1, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd3, 5'd2, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd3, 5'd3, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd3, 5'd4, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd3, 5'd5, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd3, 5'd6, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd3, 5'd7, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd4, 5'd0, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd4, 5'd1, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd4, 5'd2, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd4, 5'd3, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd4, 5'd4, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd4, 5'd5, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd4, 5'd6, 1'd0} : lccap_usb_expected = 1'b0;
  {SAS, 4'd4, 5'd7, 1'd0} : lccap_usb_expected = 1'b0;
  {PCIE, 4'd2, 5'd0, 1'd0} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd2, 5'd1, 1'd0} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd2, 5'd2, 1'd0} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd2, 5'd3, 1'd0} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd2, 5'd4, 1'd0} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd2, 5'd5, 1'd0} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd2, 5'd6, 1'd0} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd2, 5'd7, 1'd0} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd3, 5'd0, 1'd0} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd3, 5'd1, 1'd0} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd3, 5'd2, 1'd0} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd3, 5'd3, 1'd0} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd3, 5'd4, 1'd0} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd3, 5'd5, 1'd0} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd3, 5'd6, 1'd0} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd3, 5'd7, 1'd0} : lccap_usb_expected = 1'b1;
  {USB, 4'd1, 5'd0, 1'd1} : lccap_usb_expected = 1'b0;
  {USB, 4'd1, 5'd1, 1'd1} : lccap_usb_expected = 1'b0;
  {USB, 4'd1, 5'd2, 1'd1} : lccap_usb_expected = 1'b0;
  {USB, 4'd1, 5'd3, 1'd1} : lccap_usb_expected = 1'b0;
  {USB, 4'd1, 5'd4, 1'd1} : lccap_usb_expected = 1'b0;
  {USB, 4'd1, 5'd5, 1'd1} : lccap_usb_expected = 1'b0;
  {USB, 4'd1, 5'd6, 1'd1} : lccap_usb_expected = 1'b0;
  {USB, 4'd1, 5'd7, 1'd1} : lccap_usb_expected = 1'b0;
  {USB, 4'd2, 5'd0, 1'd1} : lccap_usb_expected = 1'b0;
  {USB, 4'd2, 5'd1, 1'd1} : lccap_usb_expected = 1'b0;
  {USB, 4'd2, 5'd2, 1'd1} : lccap_usb_expected = 1'b0;
  {USB, 4'd2, 5'd3, 1'd1} : lccap_usb_expected = 1'b0;
  {USB, 4'd2, 5'd4, 1'd1} : lccap_usb_expected = 1'b0;
  {USB, 4'd2, 5'd5, 1'd1} : lccap_usb_expected = 1'b0;
  {USB, 4'd2, 5'd6, 1'd1} : lccap_usb_expected = 1'b0;
  {USB, 4'd2, 5'd7, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd0, 5'd0, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd0, 5'd1, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd0, 5'd2, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd0, 5'd3, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd0, 5'd4, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd0, 5'd5, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd0, 5'd6, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd0, 5'd7, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd1, 5'd0, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd1, 5'd1, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd1, 5'd2, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd1, 5'd3, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd1, 5'd4, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd1, 5'd5, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd1, 5'd6, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd1, 5'd7, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd2, 5'd0, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd2, 5'd1, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd2, 5'd2, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd2, 5'd3, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd2, 5'd4, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd2, 5'd5, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd2, 5'd6, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd2, 5'd7, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd3, 5'd0, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd3, 5'd1, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd3, 5'd2, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd3, 5'd3, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd3, 5'd4, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd3, 5'd5, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd3, 5'd6, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd3, 5'd7, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd4, 5'd0, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd4, 5'd1, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd4, 5'd2, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd4, 5'd3, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd4, 5'd4, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd4, 5'd5, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd4, 5'd6, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd4, 5'd7, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd5, 5'd0, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd5, 5'd1, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd5, 5'd2, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd5, 5'd3, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd5, 5'd4, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd5, 5'd5, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd5, 5'd6, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd5, 5'd7, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd6, 5'd0, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd6, 5'd1, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd6, 5'd2, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd6, 5'd3, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd6, 5'd4, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd6, 5'd5, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd6, 5'd6, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd6, 5'd7, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd7, 5'd0, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd7, 5'd1, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd7, 5'd2, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd7, 5'd3, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd7, 5'd4, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd7, 5'd5, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd7, 5'd6, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd7, 5'd7, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd8, 5'd0, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd8, 5'd1, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd8, 5'd2, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd8, 5'd3, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd8, 5'd4, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd8, 5'd5, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd8, 5'd6, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd8, 5'd7, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd9, 5'd0, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd9, 5'd1, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd9, 5'd2, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd9, 5'd3, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd9, 5'd4, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd9, 5'd5, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd9, 5'd6, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd9, 5'd7, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd12, 5'd0, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd12, 5'd1, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd12, 5'd2, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd12, 5'd3, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd12, 5'd4, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd12, 5'd5, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd12, 5'd6, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd12, 5'd7, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd13, 5'd0, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd13, 5'd1, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd13, 5'd2, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd13, 5'd3, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd13, 5'd4, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd13, 5'd5, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd13, 5'd6, 1'd1} : lccap_usb_expected = 1'b0;
  {SERDES, 4'd13, 5'd7, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd0, 5'd0, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd0, 5'd1, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd0, 5'd2, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd0, 5'd3, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd0, 5'd4, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd0, 5'd5, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd0, 5'd6, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd0, 5'd7, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd1, 5'd0, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd1, 5'd1, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd1, 5'd2, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd1, 5'd3, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd1, 5'd4, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd1, 5'd5, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd1, 5'd6, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd1, 5'd7, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd2, 5'd0, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd2, 5'd1, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd2, 5'd2, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd2, 5'd3, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd2, 5'd4, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd2, 5'd5, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd2, 5'd6, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd2, 5'd7, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd3, 5'd0, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd3, 5'd1, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd3, 5'd2, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd3, 5'd3, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd3, 5'd4, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd3, 5'd5, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd3, 5'd6, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd3, 5'd7, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd4, 5'd0, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd4, 5'd1, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd4, 5'd2, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd4, 5'd3, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd4, 5'd4, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd4, 5'd5, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd4, 5'd6, 1'd1} : lccap_usb_expected = 1'b0;
  {SAS, 4'd4, 5'd7, 1'd1} : lccap_usb_expected = 1'b0;
  {PCIE, 4'd2, 5'd0, 1'd1} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd2, 5'd1, 1'd1} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd2, 5'd2, 1'd1} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd2, 5'd3, 1'd1} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd2, 5'd4, 1'd1} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd2, 5'd5, 1'd1} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd2, 5'd6, 1'd1} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd2, 5'd7, 1'd1} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd3, 5'd0, 1'd1} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd3, 5'd1, 1'd1} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd3, 5'd2, 1'd1} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd3, 5'd3, 1'd1} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd3, 5'd4, 1'd1} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd3, 5'd5, 1'd1} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd3, 5'd6, 1'd1} : lccap_usb_expected = 1'b1;
  {PCIE, 4'd3, 5'd7, 1'd1} : lccap_usb_expected = 1'b1;
default: lccap_usb_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel} )
  {USB, 4'd1, 5'd0, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd1, 5'd1, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd1, 5'd2, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd1, 5'd3, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd1, 5'd4, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd1, 5'd5, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd1, 5'd6, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd1, 5'd7, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd2, 5'd0, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd2, 5'd1, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd2, 5'd2, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd2, 5'd3, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd2, 5'd4, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd2, 5'd5, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd2, 5'd6, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd2, 5'd7, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd0, 5'd0, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd0, 5'd1, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd0, 5'd2, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd0, 5'd3, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd0, 5'd4, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd0, 5'd5, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd0, 5'd6, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd0, 5'd7, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd1, 5'd0, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd1, 5'd1, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd1, 5'd2, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd1, 5'd3, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd1, 5'd4, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd1, 5'd5, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd1, 5'd6, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd1, 5'd7, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd2, 5'd0, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd2, 5'd1, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd2, 5'd2, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd2, 5'd3, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd2, 5'd4, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd2, 5'd5, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd2, 5'd6, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd2, 5'd7, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd3, 5'd0, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd3, 5'd1, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd3, 5'd2, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd3, 5'd3, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd3, 5'd4, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd3, 5'd5, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd3, 5'd6, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd3, 5'd7, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd4, 5'd0, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd4, 5'd1, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd4, 5'd2, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd4, 5'd3, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd4, 5'd4, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd4, 5'd5, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd4, 5'd6, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd4, 5'd7, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd5, 5'd0, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd5, 5'd1, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd5, 5'd2, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd5, 5'd3, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd5, 5'd4, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd5, 5'd5, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd5, 5'd6, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd5, 5'd7, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd6, 5'd0, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd6, 5'd1, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd6, 5'd2, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd6, 5'd3, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd6, 5'd4, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd6, 5'd5, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd6, 5'd6, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd6, 5'd7, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd7, 5'd0, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd7, 5'd1, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd7, 5'd2, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd7, 5'd3, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd7, 5'd4, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd7, 5'd5, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd7, 5'd6, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd7, 5'd7, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd8, 5'd0, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd8, 5'd1, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd8, 5'd2, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd8, 5'd3, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd8, 5'd4, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd8, 5'd5, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd8, 5'd6, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd8, 5'd7, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd9, 5'd0, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd9, 5'd1, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd9, 5'd2, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd9, 5'd3, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd9, 5'd4, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd9, 5'd5, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd9, 5'd6, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd9, 5'd7, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd12, 5'd0, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd12, 5'd1, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd12, 5'd2, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd12, 5'd3, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd12, 5'd4, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd12, 5'd5, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd12, 5'd6, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd12, 5'd7, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd13, 5'd0, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd13, 5'd1, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd13, 5'd2, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd13, 5'd3, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd13, 5'd4, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd13, 5'd5, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd13, 5'd6, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd13, 5'd7, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd0, 5'd0, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd0, 5'd1, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd0, 5'd2, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd0, 5'd3, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd0, 5'd4, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd0, 5'd5, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd0, 5'd6, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd0, 5'd7, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd1, 5'd0, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd1, 5'd1, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd1, 5'd2, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd1, 5'd3, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd1, 5'd4, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd1, 5'd5, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd1, 5'd6, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd1, 5'd7, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd2, 5'd0, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd2, 5'd1, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd2, 5'd2, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd2, 5'd3, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd2, 5'd4, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd2, 5'd5, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd2, 5'd6, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd2, 5'd7, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd3, 5'd0, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd3, 5'd1, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd3, 5'd2, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd3, 5'd3, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd3, 5'd4, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd3, 5'd5, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd3, 5'd6, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd3, 5'd7, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd4, 5'd0, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd4, 5'd1, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd4, 5'd2, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd4, 5'd3, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd4, 5'd4, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd4, 5'd5, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd4, 5'd6, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd4, 5'd7, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd2, 5'd0, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd2, 5'd1, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd2, 5'd2, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd2, 5'd3, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd2, 5'd4, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd2, 5'd5, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd2, 5'd6, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd2, 5'd7, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd3, 5'd0, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd3, 5'd1, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd3, 5'd2, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd3, 5'd3, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd3, 5'd4, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd3, 5'd5, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd3, 5'd6, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd3, 5'd7, 1'd0} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd1, 5'd0, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd1, 5'd1, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd1, 5'd2, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd1, 5'd3, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd1, 5'd4, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd1, 5'd5, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd1, 5'd6, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd1, 5'd7, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd2, 5'd0, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd2, 5'd1, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd2, 5'd2, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd2, 5'd3, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd2, 5'd4, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd2, 5'd5, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd2, 5'd6, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {USB, 4'd2, 5'd7, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd0, 5'd0, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd0, 5'd1, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd0, 5'd2, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd0, 5'd3, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd0, 5'd4, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd0, 5'd5, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd0, 5'd6, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd0, 5'd7, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd1, 5'd0, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd1, 5'd1, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd1, 5'd2, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd1, 5'd3, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd1, 5'd4, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd1, 5'd5, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd1, 5'd6, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd1, 5'd7, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd2, 5'd0, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd2, 5'd1, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd2, 5'd2, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd2, 5'd3, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd2, 5'd4, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd2, 5'd5, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd2, 5'd6, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd2, 5'd7, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd3, 5'd0, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd3, 5'd1, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd3, 5'd2, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd3, 5'd3, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd3, 5'd4, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd3, 5'd5, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd3, 5'd6, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd3, 5'd7, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd4, 5'd0, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd4, 5'd1, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd4, 5'd2, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd4, 5'd3, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd4, 5'd4, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd4, 5'd5, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd4, 5'd6, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd4, 5'd7, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd5, 5'd0, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd5, 5'd1, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd5, 5'd2, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd5, 5'd3, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd5, 5'd4, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd5, 5'd5, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd5, 5'd6, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd5, 5'd7, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd6, 5'd0, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd6, 5'd1, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd6, 5'd2, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd6, 5'd3, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd6, 5'd4, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd6, 5'd5, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd6, 5'd6, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd6, 5'd7, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd7, 5'd0, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd7, 5'd1, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd7, 5'd2, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd7, 5'd3, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd7, 5'd4, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd7, 5'd5, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd7, 5'd6, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd7, 5'd7, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd8, 5'd0, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd8, 5'd1, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd8, 5'd2, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd8, 5'd3, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd8, 5'd4, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd8, 5'd5, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd8, 5'd6, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd8, 5'd7, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd9, 5'd0, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd9, 5'd1, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd9, 5'd2, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd9, 5'd3, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd9, 5'd4, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd9, 5'd5, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd9, 5'd6, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd9, 5'd7, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd12, 5'd0, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd12, 5'd1, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd12, 5'd2, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd12, 5'd3, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd12, 5'd4, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd12, 5'd5, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd12, 5'd6, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd12, 5'd7, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd13, 5'd0, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd13, 5'd1, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd13, 5'd2, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd13, 5'd3, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd13, 5'd4, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd13, 5'd5, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd13, 5'd6, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SERDES, 4'd13, 5'd7, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd0, 5'd0, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd0, 5'd1, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd0, 5'd2, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd0, 5'd3, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd0, 5'd4, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd0, 5'd5, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd0, 5'd6, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd0, 5'd7, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd1, 5'd0, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd1, 5'd1, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd1, 5'd2, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd1, 5'd3, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd1, 5'd4, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd1, 5'd5, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd1, 5'd6, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd1, 5'd7, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd2, 5'd0, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd2, 5'd1, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd2, 5'd2, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd2, 5'd3, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd2, 5'd4, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd2, 5'd5, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd2, 5'd6, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd2, 5'd7, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd3, 5'd0, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd3, 5'd1, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd3, 5'd2, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd3, 5'd3, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd3, 5'd4, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd3, 5'd5, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd3, 5'd6, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd3, 5'd7, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd4, 5'd0, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd4, 5'd1, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd4, 5'd2, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd4, 5'd3, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd4, 5'd4, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd4, 5'd5, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd4, 5'd6, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {SAS, 4'd4, 5'd7, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd2, 5'd0, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd2, 5'd1, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd2, 5'd2, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd2, 5'd3, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd2, 5'd4, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd2, 5'd5, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd2, 5'd6, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd2, 5'd7, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd3, 5'd0, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd3, 5'd1, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd3, 5'd2, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd3, 5'd3, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd3, 5'd4, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd3, 5'd5, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd3, 5'd6, 1'd1} : ssc_acc_factor_expected = 1'b0;
  {PCIE, 4'd3, 5'd7, 1'd1} : ssc_acc_factor_expected = 1'b0;
default: ssc_acc_factor_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel} )
  {USB, 4'd1, 5'd0, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {USB, 4'd1, 5'd1, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {USB, 4'd1, 5'd2, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {USB, 4'd1, 5'd3, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {USB, 4'd1, 5'd4, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {USB, 4'd1, 5'd5, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {USB, 4'd1, 5'd6, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {USB, 4'd1, 5'd7, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {USB, 4'd2, 5'd0, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {USB, 4'd2, 5'd1, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {USB, 4'd2, 5'd2, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {USB, 4'd2, 5'd3, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {USB, 4'd2, 5'd4, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {USB, 4'd2, 5'd5, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {USB, 4'd2, 5'd6, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {USB, 4'd2, 5'd7, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd0, 5'd0, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd0, 5'd1, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd0, 5'd2, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd0, 5'd3, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd0, 5'd4, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd0, 5'd5, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd0, 5'd6, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd0, 5'd7, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd1, 5'd0, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd1, 5'd1, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd1, 5'd2, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd1, 5'd3, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd1, 5'd4, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd1, 5'd5, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd1, 5'd6, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd1, 5'd7, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd2, 5'd0, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd2, 5'd1, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd2, 5'd2, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd2, 5'd3, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd2, 5'd4, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd2, 5'd5, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd2, 5'd6, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd2, 5'd7, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd3, 5'd0, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd3, 5'd1, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd3, 5'd2, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd3, 5'd3, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd3, 5'd4, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd3, 5'd5, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd3, 5'd6, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd3, 5'd7, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd4, 5'd0, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd4, 5'd1, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd4, 5'd2, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd4, 5'd3, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd4, 5'd4, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd4, 5'd5, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd4, 5'd6, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd4, 5'd7, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd5, 5'd0, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd5, 5'd1, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd5, 5'd2, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd5, 5'd3, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd5, 5'd4, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd5, 5'd5, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd5, 5'd6, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd5, 5'd7, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd6, 5'd0, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd6, 5'd1, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd6, 5'd2, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd6, 5'd3, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd6, 5'd4, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd6, 5'd5, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd6, 5'd6, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd6, 5'd7, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd7, 5'd0, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd7, 5'd1, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd7, 5'd2, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd7, 5'd3, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd7, 5'd4, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd7, 5'd5, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd7, 5'd6, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd7, 5'd7, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd8, 5'd0, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd8, 5'd1, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd8, 5'd2, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd8, 5'd3, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd8, 5'd4, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd8, 5'd5, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd8, 5'd6, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd8, 5'd7, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd9, 5'd0, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd9, 5'd1, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd9, 5'd2, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd9, 5'd3, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd9, 5'd4, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd9, 5'd5, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd9, 5'd6, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd9, 5'd7, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd12, 5'd0, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd12, 5'd1, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd12, 5'd2, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd12, 5'd3, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd12, 5'd4, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd12, 5'd5, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd12, 5'd6, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd12, 5'd7, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd13, 5'd0, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd13, 5'd1, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd13, 5'd2, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd13, 5'd3, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd13, 5'd4, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd13, 5'd5, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd13, 5'd6, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SERDES, 4'd13, 5'd7, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd0, 5'd0, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd0, 5'd1, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd0, 5'd2, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd0, 5'd3, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd0, 5'd4, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd0, 5'd5, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd0, 5'd6, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd0, 5'd7, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd1, 5'd0, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd1, 5'd1, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd1, 5'd2, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd1, 5'd3, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd1, 5'd4, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd1, 5'd5, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd1, 5'd6, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd1, 5'd7, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd2, 5'd0, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd2, 5'd1, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd2, 5'd2, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd2, 5'd3, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd2, 5'd4, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd2, 5'd5, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd2, 5'd6, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd2, 5'd7, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd3, 5'd0, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd3, 5'd1, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd3, 5'd2, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd3, 5'd3, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd3, 5'd4, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd3, 5'd5, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd3, 5'd6, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd3, 5'd7, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd4, 5'd0, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd4, 5'd1, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd4, 5'd2, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd4, 5'd3, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd4, 5'd4, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd4, 5'd5, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd4, 5'd6, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {SAS, 4'd4, 5'd7, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {PCIE, 4'd2, 5'd0, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {PCIE, 4'd2, 5'd1, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {PCIE, 4'd2, 5'd2, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {PCIE, 4'd2, 5'd3, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {PCIE, 4'd2, 5'd4, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {PCIE, 4'd2, 5'd5, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {PCIE, 4'd2, 5'd6, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {PCIE, 4'd2, 5'd7, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {PCIE, 4'd3, 5'd0, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {PCIE, 4'd3, 5'd1, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {PCIE, 4'd3, 5'd2, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {PCIE, 4'd3, 5'd3, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {PCIE, 4'd3, 5'd4, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {PCIE, 4'd3, 5'd5, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {PCIE, 4'd3, 5'd6, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {PCIE, 4'd3, 5'd7, 1'd0} : ssc_step_125ppm_expected = 4'b0000;
  {USB, 4'd1, 5'd0, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {USB, 4'd1, 5'd1, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {USB, 4'd1, 5'd2, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {USB, 4'd1, 5'd3, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {USB, 4'd1, 5'd4, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {USB, 4'd1, 5'd5, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {USB, 4'd1, 5'd6, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {USB, 4'd1, 5'd7, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {USB, 4'd2, 5'd0, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {USB, 4'd2, 5'd1, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {USB, 4'd2, 5'd2, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {USB, 4'd2, 5'd3, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {USB, 4'd2, 5'd4, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {USB, 4'd2, 5'd5, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {USB, 4'd2, 5'd6, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {USB, 4'd2, 5'd7, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd0, 5'd0, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd0, 5'd1, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd0, 5'd2, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd0, 5'd3, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd0, 5'd4, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd0, 5'd5, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd0, 5'd6, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd0, 5'd7, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd1, 5'd0, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd1, 5'd1, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd1, 5'd2, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd1, 5'd3, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd1, 5'd4, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd1, 5'd5, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd1, 5'd6, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd1, 5'd7, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd2, 5'd0, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd2, 5'd1, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd2, 5'd2, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd2, 5'd3, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd2, 5'd4, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd2, 5'd5, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd2, 5'd6, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd2, 5'd7, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd3, 5'd0, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd3, 5'd1, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd3, 5'd2, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd3, 5'd3, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd3, 5'd4, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd3, 5'd5, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd3, 5'd6, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd3, 5'd7, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd4, 5'd0, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd4, 5'd1, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd4, 5'd2, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd4, 5'd3, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd4, 5'd4, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd4, 5'd5, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd4, 5'd6, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd4, 5'd7, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd5, 5'd0, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd5, 5'd1, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd5, 5'd2, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd5, 5'd3, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd5, 5'd4, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd5, 5'd5, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd5, 5'd6, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd5, 5'd7, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd6, 5'd0, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd6, 5'd1, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd6, 5'd2, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd6, 5'd3, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd6, 5'd4, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd6, 5'd5, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd6, 5'd6, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd6, 5'd7, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd7, 5'd0, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd7, 5'd1, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd7, 5'd2, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd7, 5'd3, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd7, 5'd4, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd7, 5'd5, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd7, 5'd6, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd7, 5'd7, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd8, 5'd0, 1'd1} : ssc_step_125ppm_expected = 4'b0010;
  {SERDES, 4'd8, 5'd1, 1'd1} : ssc_step_125ppm_expected = 4'b0010;
  {SERDES, 4'd8, 5'd2, 1'd1} : ssc_step_125ppm_expected = 4'b0010;
  {SERDES, 4'd8, 5'd3, 1'd1} : ssc_step_125ppm_expected = 4'b0010;
  {SERDES, 4'd8, 5'd4, 1'd1} : ssc_step_125ppm_expected = 4'b0010;
  {SERDES, 4'd8, 5'd5, 1'd1} : ssc_step_125ppm_expected = 4'b0010;
  {SERDES, 4'd8, 5'd6, 1'd1} : ssc_step_125ppm_expected = 4'b0010;
  {SERDES, 4'd8, 5'd7, 1'd1} : ssc_step_125ppm_expected = 4'b0010;
  {SERDES, 4'd9, 5'd0, 1'd1} : ssc_step_125ppm_expected = 4'b0010;
  {SERDES, 4'd9, 5'd1, 1'd1} : ssc_step_125ppm_expected = 4'b0010;
  {SERDES, 4'd9, 5'd2, 1'd1} : ssc_step_125ppm_expected = 4'b0010;
  {SERDES, 4'd9, 5'd3, 1'd1} : ssc_step_125ppm_expected = 4'b0010;
  {SERDES, 4'd9, 5'd4, 1'd1} : ssc_step_125ppm_expected = 4'b0010;
  {SERDES, 4'd9, 5'd5, 1'd1} : ssc_step_125ppm_expected = 4'b0010;
  {SERDES, 4'd9, 5'd6, 1'd1} : ssc_step_125ppm_expected = 4'b0010;
  {SERDES, 4'd9, 5'd7, 1'd1} : ssc_step_125ppm_expected = 4'b0010;
  {SERDES, 4'd12, 5'd0, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd12, 5'd1, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd12, 5'd2, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd12, 5'd3, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd12, 5'd4, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd12, 5'd5, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd12, 5'd6, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd12, 5'd7, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd13, 5'd0, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd13, 5'd1, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd13, 5'd2, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd13, 5'd3, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd13, 5'd4, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd13, 5'd5, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd13, 5'd6, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SERDES, 4'd13, 5'd7, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd0, 5'd0, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd0, 5'd1, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd0, 5'd2, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd0, 5'd3, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd0, 5'd4, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd0, 5'd5, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd0, 5'd6, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd0, 5'd7, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd1, 5'd0, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd1, 5'd1, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd1, 5'd2, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd1, 5'd3, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd1, 5'd4, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd1, 5'd5, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd1, 5'd6, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd1, 5'd7, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd2, 5'd0, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd2, 5'd1, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd2, 5'd2, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd2, 5'd3, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd2, 5'd4, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd2, 5'd5, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd2, 5'd6, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd2, 5'd7, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd3, 5'd0, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd3, 5'd1, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd3, 5'd2, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd3, 5'd3, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd3, 5'd4, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd3, 5'd5, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd3, 5'd6, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd3, 5'd7, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd4, 5'd0, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd4, 5'd1, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd4, 5'd2, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd4, 5'd3, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd4, 5'd4, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd4, 5'd5, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd4, 5'd6, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {SAS, 4'd4, 5'd7, 1'd1} : ssc_step_125ppm_expected = 4'b0011;
  {PCIE, 4'd2, 5'd0, 1'd1} : ssc_step_125ppm_expected = 4'b0100;
  {PCIE, 4'd2, 5'd1, 1'd1} : ssc_step_125ppm_expected = 4'b0100;
  {PCIE, 4'd2, 5'd2, 1'd1} : ssc_step_125ppm_expected = 4'b0100;
  {PCIE, 4'd2, 5'd3, 1'd1} : ssc_step_125ppm_expected = 4'b0100;
  {PCIE, 4'd2, 5'd4, 1'd1} : ssc_step_125ppm_expected = 4'b0100;
  {PCIE, 4'd2, 5'd5, 1'd1} : ssc_step_125ppm_expected = 4'b0100;
  {PCIE, 4'd2, 5'd6, 1'd1} : ssc_step_125ppm_expected = 4'b0100;
  {PCIE, 4'd2, 5'd7, 1'd1} : ssc_step_125ppm_expected = 4'b0100;
  {PCIE, 4'd3, 5'd0, 1'd1} : ssc_step_125ppm_expected = 4'b0100;
  {PCIE, 4'd3, 5'd1, 1'd1} : ssc_step_125ppm_expected = 4'b0100;
  {PCIE, 4'd3, 5'd2, 1'd1} : ssc_step_125ppm_expected = 4'b0100;
  {PCIE, 4'd3, 5'd3, 1'd1} : ssc_step_125ppm_expected = 4'b0100;
  {PCIE, 4'd3, 5'd4, 1'd1} : ssc_step_125ppm_expected = 4'b0100;
  {PCIE, 4'd3, 5'd5, 1'd1} : ssc_step_125ppm_expected = 4'b0100;
  {PCIE, 4'd3, 5'd6, 1'd1} : ssc_step_125ppm_expected = 4'b0100;
  {PCIE, 4'd3, 5'd7, 1'd1} : ssc_step_125ppm_expected = 4'b0100;
default: ssc_step_125ppm_expected = 4'bzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel[4:0], reg_fbck_sel} )
  {USB, 4'd1, 5'd0, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd1, 5'd1, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd1, 5'd2, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd1, 5'd3, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd1, 5'd4, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd1, 5'd5, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd1, 5'd6, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd1, 5'd7, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd2, 5'd0, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd2, 5'd1, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd2, 5'd2, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd2, 5'd3, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd2, 5'd4, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd2, 5'd5, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd2, 5'd6, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd2, 5'd7, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd0, 5'd0, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd0, 5'd1, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd0, 5'd2, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd0, 5'd3, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd0, 5'd4, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd0, 5'd5, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd0, 5'd6, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd0, 5'd7, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd1, 5'd0, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd1, 5'd1, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd1, 5'd2, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd1, 5'd3, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd1, 5'd4, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd1, 5'd5, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd1, 5'd6, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd1, 5'd7, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd2, 5'd0, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd2, 5'd1, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd2, 5'd2, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd2, 5'd3, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd2, 5'd4, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd2, 5'd5, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd2, 5'd6, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd2, 5'd7, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd3, 5'd0, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd3, 5'd1, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd3, 5'd2, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd3, 5'd3, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd3, 5'd4, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd3, 5'd5, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd3, 5'd6, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd3, 5'd7, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd4, 5'd0, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd4, 5'd1, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd4, 5'd2, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd4, 5'd3, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd4, 5'd4, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd4, 5'd5, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd4, 5'd6, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd4, 5'd7, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd5, 5'd0, 1'd0} : ssc_m_expected = 13'b0101111001101;
  {SERDES, 4'd5, 5'd1, 1'd0} : ssc_m_expected = 13'b0101111001101;
  {SERDES, 4'd5, 5'd2, 1'd0} : ssc_m_expected = 13'b0101111001101;
  {SERDES, 4'd5, 5'd3, 1'd0} : ssc_m_expected = 13'b0101111001101;
  {SERDES, 4'd5, 5'd4, 1'd0} : ssc_m_expected = 13'b0101111001101;
  {SERDES, 4'd5, 5'd5, 1'd0} : ssc_m_expected = 13'b0101111001101;
  {SERDES, 4'd5, 5'd6, 1'd0} : ssc_m_expected = 13'b0101111001101;
  {SERDES, 4'd5, 5'd7, 1'd0} : ssc_m_expected = 13'b0101111001101;
  {SERDES, 4'd6, 5'd0, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd6, 5'd1, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd6, 5'd2, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd6, 5'd3, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd6, 5'd4, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd6, 5'd5, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd6, 5'd6, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd6, 5'd7, 1'd0} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd7, 5'd0, 1'd0} : ssc_m_expected = 13'b0110001111011;
  {SERDES, 4'd7, 5'd1, 1'd0} : ssc_m_expected = 13'b0110001111011;
  {SERDES, 4'd7, 5'd2, 1'd0} : ssc_m_expected = 13'b0110001111011;
  {SERDES, 4'd7, 5'd3, 1'd0} : ssc_m_expected = 13'b0110001111011;
  {SERDES, 4'd7, 5'd4, 1'd0} : ssc_m_expected = 13'b0110001111011;
  {SERDES, 4'd7, 5'd5, 1'd0} : ssc_m_expected = 13'b0110001111011;
  {SERDES, 4'd7, 5'd6, 1'd0} : ssc_m_expected = 13'b0110001111011;
  {SERDES, 4'd7, 5'd7, 1'd0} : ssc_m_expected = 13'b0110001111011;
  {SERDES, 4'd8, 5'd0, 1'd0} : ssc_m_expected = 13'b0110101010001;
  {SERDES, 4'd8, 5'd1, 1'd0} : ssc_m_expected = 13'b0110101010001;
  {SERDES, 4'd8, 5'd2, 1'd0} : ssc_m_expected = 13'b0110101010001;
  {SERDES, 4'd8, 5'd3, 1'd0} : ssc_m_expected = 13'b0110101010001;
  {SERDES, 4'd8, 5'd4, 1'd0} : ssc_m_expected = 13'b0110101010001;
  {SERDES, 4'd8, 5'd5, 1'd0} : ssc_m_expected = 13'b0110101010001;
  {SERDES, 4'd8, 5'd6, 1'd0} : ssc_m_expected = 13'b0110101010001;
  {SERDES, 4'd8, 5'd7, 1'd0} : ssc_m_expected = 13'b0110101010001;
  {SERDES, 4'd9, 5'd0, 1'd0} : ssc_m_expected = 13'b0110110011101;
  {SERDES, 4'd9, 5'd1, 1'd0} : ssc_m_expected = 13'b0110110011101;
  {SERDES, 4'd9, 5'd2, 1'd0} : ssc_m_expected = 13'b0110110011101;
  {SERDES, 4'd9, 5'd3, 1'd0} : ssc_m_expected = 13'b0110110011101;
  {SERDES, 4'd9, 5'd4, 1'd0} : ssc_m_expected = 13'b0110110011101;
  {SERDES, 4'd9, 5'd5, 1'd0} : ssc_m_expected = 13'b0110110011101;
  {SERDES, 4'd9, 5'd6, 1'd0} : ssc_m_expected = 13'b0110110011101;
  {SERDES, 4'd9, 5'd7, 1'd0} : ssc_m_expected = 13'b0110110011101;
  {SERDES, 4'd12, 5'd0, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd12, 5'd1, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd12, 5'd2, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd12, 5'd3, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd12, 5'd4, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd12, 5'd5, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd12, 5'd6, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd12, 5'd7, 1'd0} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd13, 5'd0, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd13, 5'd1, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd13, 5'd2, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd13, 5'd3, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd13, 5'd4, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd13, 5'd5, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd13, 5'd6, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd13, 5'd7, 1'd0} : ssc_m_expected = 13'b0100111111011;
  {SAS, 4'd0, 5'd0, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd0, 5'd1, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd0, 5'd2, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd0, 5'd3, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd0, 5'd4, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd0, 5'd5, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd0, 5'd6, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd0, 5'd7, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd1, 5'd0, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd1, 5'd1, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd1, 5'd2, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd1, 5'd3, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd1, 5'd4, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd1, 5'd5, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd1, 5'd6, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd1, 5'd7, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd2, 5'd0, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd2, 5'd1, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd2, 5'd2, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd2, 5'd3, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd2, 5'd4, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd2, 5'd5, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd2, 5'd6, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd2, 5'd7, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd3, 5'd0, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd3, 5'd1, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd3, 5'd2, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd3, 5'd3, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd3, 5'd4, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd3, 5'd5, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd3, 5'd6, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd3, 5'd7, 1'd0} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd4, 5'd0, 1'd0} : ssc_m_expected = 13'b0101011100101;
  {SAS, 4'd4, 5'd1, 1'd0} : ssc_m_expected = 13'b0101011100101;
  {SAS, 4'd4, 5'd2, 1'd0} : ssc_m_expected = 13'b0101011100101;
  {SAS, 4'd4, 5'd3, 1'd0} : ssc_m_expected = 13'b0101011100101;
  {SAS, 4'd4, 5'd4, 1'd0} : ssc_m_expected = 13'b0101011100101;
  {SAS, 4'd4, 5'd5, 1'd0} : ssc_m_expected = 13'b0101011100101;
  {SAS, 4'd4, 5'd6, 1'd0} : ssc_m_expected = 13'b0101011100101;
  {SAS, 4'd4, 5'd7, 1'd0} : ssc_m_expected = 13'b0101011100101;
  {PCIE, 4'd2, 5'd0, 1'd0} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd2, 5'd1, 1'd0} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd2, 5'd2, 1'd0} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd2, 5'd3, 1'd0} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd2, 5'd4, 1'd0} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd2, 5'd5, 1'd0} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd2, 5'd6, 1'd0} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd2, 5'd7, 1'd0} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd3, 5'd0, 1'd0} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd3, 5'd1, 1'd0} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd3, 5'd2, 1'd0} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd3, 5'd3, 1'd0} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd3, 5'd4, 1'd0} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd3, 5'd5, 1'd0} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd3, 5'd6, 1'd0} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd3, 5'd7, 1'd0} : ssc_m_expected = 13'b0011110111111;
  {USB, 4'd1, 5'd0, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd1, 5'd1, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd1, 5'd2, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd1, 5'd3, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd1, 5'd4, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd1, 5'd5, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd1, 5'd6, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd1, 5'd7, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd2, 5'd0, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd2, 5'd1, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd2, 5'd2, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd2, 5'd3, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd2, 5'd4, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd2, 5'd5, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd2, 5'd6, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {USB, 4'd2, 5'd7, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd0, 5'd0, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd0, 5'd1, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd0, 5'd2, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd0, 5'd3, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd0, 5'd4, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd0, 5'd5, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd0, 5'd6, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd0, 5'd7, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd1, 5'd0, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd1, 5'd1, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd1, 5'd2, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd1, 5'd3, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd1, 5'd4, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd1, 5'd5, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd1, 5'd6, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd1, 5'd7, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd2, 5'd0, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd2, 5'd1, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd2, 5'd2, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd2, 5'd3, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd2, 5'd4, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd2, 5'd5, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd2, 5'd6, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd2, 5'd7, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd3, 5'd0, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd3, 5'd1, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd3, 5'd2, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd3, 5'd3, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd3, 5'd4, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd3, 5'd5, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd3, 5'd6, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd3, 5'd7, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd4, 5'd0, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd4, 5'd1, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd4, 5'd2, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd4, 5'd3, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd4, 5'd4, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd4, 5'd5, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd4, 5'd6, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd4, 5'd7, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd5, 5'd0, 1'd1} : ssc_m_expected = 13'b0101111001101;
  {SERDES, 4'd5, 5'd1, 1'd1} : ssc_m_expected = 13'b0101111001101;
  {SERDES, 4'd5, 5'd2, 1'd1} : ssc_m_expected = 13'b0101111001101;
  {SERDES, 4'd5, 5'd3, 1'd1} : ssc_m_expected = 13'b0101111001101;
  {SERDES, 4'd5, 5'd4, 1'd1} : ssc_m_expected = 13'b0101111001101;
  {SERDES, 4'd5, 5'd5, 1'd1} : ssc_m_expected = 13'b0101111001101;
  {SERDES, 4'd5, 5'd6, 1'd1} : ssc_m_expected = 13'b0101111001101;
  {SERDES, 4'd5, 5'd7, 1'd1} : ssc_m_expected = 13'b0101111001101;
  {SERDES, 4'd6, 5'd0, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd6, 5'd1, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd6, 5'd2, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd6, 5'd3, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd6, 5'd4, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd6, 5'd5, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd6, 5'd6, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd6, 5'd7, 1'd1} : ssc_m_expected = 13'b0110000011011;
  {SERDES, 4'd7, 5'd0, 1'd1} : ssc_m_expected = 13'b0110001111011;
  {SERDES, 4'd7, 5'd1, 1'd1} : ssc_m_expected = 13'b0110001111011;
  {SERDES, 4'd7, 5'd2, 1'd1} : ssc_m_expected = 13'b0110001111011;
  {SERDES, 4'd7, 5'd3, 1'd1} : ssc_m_expected = 13'b0110001111011;
  {SERDES, 4'd7, 5'd4, 1'd1} : ssc_m_expected = 13'b0110001111011;
  {SERDES, 4'd7, 5'd5, 1'd1} : ssc_m_expected = 13'b0110001111011;
  {SERDES, 4'd7, 5'd6, 1'd1} : ssc_m_expected = 13'b0110001111011;
  {SERDES, 4'd7, 5'd7, 1'd1} : ssc_m_expected = 13'b0110001111011;
  {SERDES, 4'd8, 5'd0, 1'd1} : ssc_m_expected = 13'b0110101010001;
  {SERDES, 4'd8, 5'd1, 1'd1} : ssc_m_expected = 13'b0110101010001;
  {SERDES, 4'd8, 5'd2, 1'd1} : ssc_m_expected = 13'b0110101010001;
  {SERDES, 4'd8, 5'd3, 1'd1} : ssc_m_expected = 13'b0110101010001;
  {SERDES, 4'd8, 5'd4, 1'd1} : ssc_m_expected = 13'b0110101010001;
  {SERDES, 4'd8, 5'd5, 1'd1} : ssc_m_expected = 13'b0110101010001;
  {SERDES, 4'd8, 5'd6, 1'd1} : ssc_m_expected = 13'b0110101010001;
  {SERDES, 4'd8, 5'd7, 1'd1} : ssc_m_expected = 13'b0110101010001;
  {SERDES, 4'd9, 5'd0, 1'd1} : ssc_m_expected = 13'b0110110011101;
  {SERDES, 4'd9, 5'd1, 1'd1} : ssc_m_expected = 13'b0110110011101;
  {SERDES, 4'd9, 5'd2, 1'd1} : ssc_m_expected = 13'b0110110011101;
  {SERDES, 4'd9, 5'd3, 1'd1} : ssc_m_expected = 13'b0110110011101;
  {SERDES, 4'd9, 5'd4, 1'd1} : ssc_m_expected = 13'b0110110011101;
  {SERDES, 4'd9, 5'd5, 1'd1} : ssc_m_expected = 13'b0110110011101;
  {SERDES, 4'd9, 5'd6, 1'd1} : ssc_m_expected = 13'b0110110011101;
  {SERDES, 4'd9, 5'd7, 1'd1} : ssc_m_expected = 13'b0110110011101;
  {SERDES, 4'd12, 5'd0, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd12, 5'd1, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd12, 5'd2, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd12, 5'd3, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd12, 5'd4, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd12, 5'd5, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd12, 5'd6, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd12, 5'd7, 1'd1} : ssc_m_expected = 13'b0100110101111;
  {SERDES, 4'd13, 5'd0, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd13, 5'd1, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd13, 5'd2, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd13, 5'd3, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd13, 5'd4, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd13, 5'd5, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd13, 5'd6, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SERDES, 4'd13, 5'd7, 1'd1} : ssc_m_expected = 13'b0100111111011;
  {SAS, 4'd0, 5'd0, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd0, 5'd1, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd0, 5'd2, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd0, 5'd3, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd0, 5'd4, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd0, 5'd5, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd0, 5'd6, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd0, 5'd7, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd1, 5'd0, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd1, 5'd1, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd1, 5'd2, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd1, 5'd3, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd1, 5'd4, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd1, 5'd5, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd1, 5'd6, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd1, 5'd7, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd2, 5'd0, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd2, 5'd1, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd2, 5'd2, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd2, 5'd3, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd2, 5'd4, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd2, 5'd5, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd2, 5'd6, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd2, 5'd7, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd3, 5'd0, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd3, 5'd1, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd3, 5'd2, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd3, 5'd3, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd3, 5'd4, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd3, 5'd5, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd3, 5'd6, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd3, 5'd7, 1'd1} : ssc_m_expected = 13'b0101110011111;
  {SAS, 4'd4, 5'd0, 1'd1} : ssc_m_expected = 13'b0101011100101;
  {SAS, 4'd4, 5'd1, 1'd1} : ssc_m_expected = 13'b0101011100101;
  {SAS, 4'd4, 5'd2, 1'd1} : ssc_m_expected = 13'b0101011100101;
  {SAS, 4'd4, 5'd3, 1'd1} : ssc_m_expected = 13'b0101011100101;
  {SAS, 4'd4, 5'd4, 1'd1} : ssc_m_expected = 13'b0101011100101;
  {SAS, 4'd4, 5'd5, 1'd1} : ssc_m_expected = 13'b0101011100101;
  {SAS, 4'd4, 5'd6, 1'd1} : ssc_m_expected = 13'b0101011100101;
  {SAS, 4'd4, 5'd7, 1'd1} : ssc_m_expected = 13'b0101011100101;
  {PCIE, 4'd2, 5'd0, 1'd1} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd2, 5'd1, 1'd1} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd2, 5'd2, 1'd1} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd2, 5'd3, 1'd1} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd2, 5'd4, 1'd1} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd2, 5'd5, 1'd1} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd2, 5'd6, 1'd1} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd2, 5'd7, 1'd1} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd3, 5'd0, 1'd1} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd3, 5'd1, 1'd1} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd3, 5'd2, 1'd1} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd3, 5'd3, 1'd1} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd3, 5'd4, 1'd1} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd3, 5'd5, 1'd1} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd3, 5'd6, 1'd1} : ssc_m_expected = 13'b0011110111111;
  {PCIE, 4'd3, 5'd7, 1'd1} : ssc_m_expected = 13'b0011110111111;
default: ssc_m_expected = 13'bzzzzzzzzzzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel} )
  {PCIE, 4'd0, 5'd0, 1'd0} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd1, 1'd0} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd2, 1'd0} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd3, 1'd0} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd4, 1'd0} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd5, 1'd0} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd6, 1'd0} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd7, 1'd0} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd0, 1'd0} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd1, 1'd0} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd2, 1'd0} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd3, 1'd0} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd4, 1'd0} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd5, 1'd0} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd6, 1'd0} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd7, 1'd0} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd0, 1'd1} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd1, 1'd1} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd2, 1'd1} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd3, 1'd1} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd4, 1'd1} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd5, 1'd1} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd6, 1'd1} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd7, 1'd1} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd0, 1'd1} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd1, 1'd1} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd2, 1'd1} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd3, 1'd1} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd4, 1'd1} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd5, 1'd1} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd6, 1'd1} : ref_clk_ring_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd7, 1'd1} : ref_clk_ring_sel_expected = 1'b1;
default: ref_clk_ring_sel_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel} )
  {PCIE, 4'd0, 5'd0, 1'd0} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd1, 1'd0} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd2, 1'd0} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd3, 1'd0} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd4, 1'd0} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd5, 1'd0} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd6, 1'd0} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd7, 1'd0} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd0, 1'd0} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd1, 1'd0} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd2, 1'd0} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd3, 1'd0} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd4, 1'd0} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd5, 1'd0} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd6, 1'd0} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd7, 1'd0} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd0, 1'd1} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd1, 1'd1} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd2, 1'd1} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd3, 1'd1} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd4, 1'd1} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd5, 1'd1} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd6, 1'd1} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd0, 5'd7, 1'd1} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd0, 1'd1} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd1, 1'd1} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd2, 1'd1} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd3, 1'd1} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd4, 1'd1} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd5, 1'd1} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd6, 1'd1} : clk1g_refclk_sel_expected = 1'b1;
  {PCIE, 4'd1, 5'd7, 1'd1} : clk1g_refclk_sel_expected = 1'b1;
default: clk1g_refclk_sel_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel} )
  {PCIE, 4'd0, 5'd0, 1'd0} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd0, 5'd1, 1'd0} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd0, 5'd2, 1'd0} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd0, 5'd3, 1'd0} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd0, 5'd4, 1'd0} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd0, 5'd5, 1'd0} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd0, 5'd6, 1'd0} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd0, 5'd7, 1'd0} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd1, 5'd0, 1'd0} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd1, 5'd1, 1'd0} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd1, 5'd2, 1'd0} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd1, 5'd3, 1'd0} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd1, 5'd4, 1'd0} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd1, 5'd5, 1'd0} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd1, 5'd6, 1'd0} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd1, 5'd7, 1'd0} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd0, 5'd0, 1'd1} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd0, 5'd1, 1'd1} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd0, 5'd2, 1'd1} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd0, 5'd3, 1'd1} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd0, 5'd4, 1'd1} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd0, 5'd5, 1'd1} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd0, 5'd6, 1'd1} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd0, 5'd7, 1'd1} : pll_refdiv_ring_expected = 4'b0010;
  {PCIE, 4'd1, 5'd0, 1'd1} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd1, 5'd1, 1'd1} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd1, 5'd2, 1'd1} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd1, 5'd3, 1'd1} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd1, 5'd4, 1'd1} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd1, 5'd5, 1'd1} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd1, 5'd6, 1'd1} : pll_refdiv_ring_expected = 4'b0001;
  {PCIE, 4'd1, 5'd7, 1'd1} : pll_refdiv_ring_expected = 4'b0010;
default: pll_refdiv_ring_expected = 4'bzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel} )
  {PCIE, 4'd0, 5'd0, 1'd0} : pll_fbdiv_ring_expected = 10'b0110010000;
  {PCIE, 4'd0, 5'd1, 1'd0} : pll_fbdiv_ring_expected = 10'b0101001101;
  {PCIE, 4'd0, 5'd2, 1'd0} : pll_fbdiv_ring_expected = 10'b0011111010;
  {PCIE, 4'd0, 5'd3, 1'd0} : pll_fbdiv_ring_expected = 10'b0011001000;
  {PCIE, 4'd0, 5'd4, 1'd0} : pll_fbdiv_ring_expected = 10'b0010100000;
  {PCIE, 4'd0, 5'd5, 1'd0} : pll_fbdiv_ring_expected = 10'b0001100100;
  {PCIE, 4'd0, 5'd6, 1'd0} : pll_fbdiv_ring_expected = 10'b0001010000;
  {PCIE, 4'd0, 5'd7, 1'd0} : pll_fbdiv_ring_expected = 10'b0001000000;
  {PCIE, 4'd1, 5'd0, 1'd0} : pll_fbdiv_ring_expected = 10'b0110010000;
  {PCIE, 4'd1, 5'd1, 1'd0} : pll_fbdiv_ring_expected = 10'b0101001101;
  {PCIE, 4'd1, 5'd2, 1'd0} : pll_fbdiv_ring_expected = 10'b0011111010;
  {PCIE, 4'd1, 5'd3, 1'd0} : pll_fbdiv_ring_expected = 10'b0011001000;
  {PCIE, 4'd1, 5'd4, 1'd0} : pll_fbdiv_ring_expected = 10'b0010100000;
  {PCIE, 4'd1, 5'd5, 1'd0} : pll_fbdiv_ring_expected = 10'b0001100100;
  {PCIE, 4'd1, 5'd6, 1'd0} : pll_fbdiv_ring_expected = 10'b0001010000;
  {PCIE, 4'd1, 5'd7, 1'd0} : pll_fbdiv_ring_expected = 10'b0001000000;
  {PCIE, 4'd0, 5'd0, 1'd1} : pll_fbdiv_ring_expected = 10'b0001100100;
  {PCIE, 4'd0, 5'd1, 1'd1} : pll_fbdiv_ring_expected = 10'b0001010011;
  {PCIE, 4'd0, 5'd2, 1'd1} : pll_fbdiv_ring_expected = 10'b0000111110;
  {PCIE, 4'd0, 5'd3, 1'd1} : pll_fbdiv_ring_expected = 10'b0000110010;
  {PCIE, 4'd0, 5'd4, 1'd1} : pll_fbdiv_ring_expected = 10'b0000101000;
  {PCIE, 4'd0, 5'd5, 1'd1} : pll_fbdiv_ring_expected = 10'b0000011001;
  {PCIE, 4'd0, 5'd6, 1'd1} : pll_fbdiv_ring_expected = 10'b0000010100;
  {PCIE, 4'd0, 5'd7, 1'd1} : pll_fbdiv_ring_expected = 10'b0000100000;
  {PCIE, 4'd1, 5'd0, 1'd1} : pll_fbdiv_ring_expected = 10'b0001100100;
  {PCIE, 4'd1, 5'd1, 1'd1} : pll_fbdiv_ring_expected = 10'b0001010011;
  {PCIE, 4'd1, 5'd2, 1'd1} : pll_fbdiv_ring_expected = 10'b0000111110;
  {PCIE, 4'd1, 5'd3, 1'd1} : pll_fbdiv_ring_expected = 10'b0000110010;
  {PCIE, 4'd1, 5'd4, 1'd1} : pll_fbdiv_ring_expected = 10'b0000101000;
  {PCIE, 4'd1, 5'd5, 1'd1} : pll_fbdiv_ring_expected = 10'b0000011001;
  {PCIE, 4'd1, 5'd6, 1'd1} : pll_fbdiv_ring_expected = 10'b0000010100;
  {PCIE, 4'd1, 5'd7, 1'd1} : pll_fbdiv_ring_expected = 10'b0000100000;
default: pll_fbdiv_ring_expected = 10'bzzzzzzzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel} )
  {PCIE, 4'd0, 5'd0, 1'd0} : pll_fbdiv_ring_fbck_expected = 10'b0110010000;
  {PCIE, 4'd0, 5'd1, 1'd0} : pll_fbdiv_ring_fbck_expected = 10'b0101001101;
  {PCIE, 4'd0, 5'd2, 1'd0} : pll_fbdiv_ring_fbck_expected = 10'b0011111010;
  {PCIE, 4'd0, 5'd3, 1'd0} : pll_fbdiv_ring_fbck_expected = 10'b0011001000;
  {PCIE, 4'd0, 5'd4, 1'd0} : pll_fbdiv_ring_fbck_expected = 10'b0010100000;
  {PCIE, 4'd0, 5'd5, 1'd0} : pll_fbdiv_ring_fbck_expected = 10'b0001100100;
  {PCIE, 4'd0, 5'd6, 1'd0} : pll_fbdiv_ring_fbck_expected = 10'b0001010000;
  {PCIE, 4'd0, 5'd7, 1'd0} : pll_fbdiv_ring_fbck_expected = 10'b0001000000;
  {PCIE, 4'd1, 5'd0, 1'd0} : pll_fbdiv_ring_fbck_expected = 10'b0110010000;
  {PCIE, 4'd1, 5'd1, 1'd0} : pll_fbdiv_ring_fbck_expected = 10'b0101001101;
  {PCIE, 4'd1, 5'd2, 1'd0} : pll_fbdiv_ring_fbck_expected = 10'b0011111010;
  {PCIE, 4'd1, 5'd3, 1'd0} : pll_fbdiv_ring_fbck_expected = 10'b0011001000;
  {PCIE, 4'd1, 5'd4, 1'd0} : pll_fbdiv_ring_fbck_expected = 10'b0010100000;
  {PCIE, 4'd1, 5'd5, 1'd0} : pll_fbdiv_ring_fbck_expected = 10'b0001100100;
  {PCIE, 4'd1, 5'd6, 1'd0} : pll_fbdiv_ring_fbck_expected = 10'b0001010000;
  {PCIE, 4'd1, 5'd7, 1'd0} : pll_fbdiv_ring_fbck_expected = 10'b0001000000;
  {PCIE, 4'd0, 5'd0, 1'd1} : pll_fbdiv_ring_fbck_expected = 10'b0001100100;
  {PCIE, 4'd0, 5'd1, 1'd1} : pll_fbdiv_ring_fbck_expected = 10'b0001010011;
  {PCIE, 4'd0, 5'd2, 1'd1} : pll_fbdiv_ring_fbck_expected = 10'b0000111110;
  {PCIE, 4'd0, 5'd3, 1'd1} : pll_fbdiv_ring_fbck_expected = 10'b0000110010;
  {PCIE, 4'd0, 5'd4, 1'd1} : pll_fbdiv_ring_fbck_expected = 10'b0000101000;
  {PCIE, 4'd0, 5'd5, 1'd1} : pll_fbdiv_ring_fbck_expected = 10'b0000011001;
  {PCIE, 4'd0, 5'd6, 1'd1} : pll_fbdiv_ring_fbck_expected = 10'b0000010100;
  {PCIE, 4'd0, 5'd7, 1'd1} : pll_fbdiv_ring_fbck_expected = 10'b0000100000;
  {PCIE, 4'd1, 5'd0, 1'd1} : pll_fbdiv_ring_fbck_expected = 10'b0001100100;
  {PCIE, 4'd1, 5'd1, 1'd1} : pll_fbdiv_ring_fbck_expected = 10'b0001010011;
  {PCIE, 4'd1, 5'd2, 1'd1} : pll_fbdiv_ring_fbck_expected = 10'b0000111110;
  {PCIE, 4'd1, 5'd3, 1'd1} : pll_fbdiv_ring_fbck_expected = 10'b0000110010;
  {PCIE, 4'd1, 5'd4, 1'd1} : pll_fbdiv_ring_fbck_expected = 10'b0000101000;
  {PCIE, 4'd1, 5'd5, 1'd1} : pll_fbdiv_ring_fbck_expected = 10'b0000011001;
  {PCIE, 4'd1, 5'd6, 1'd1} : pll_fbdiv_ring_fbck_expected = 10'b0000010100;
  {PCIE, 4'd1, 5'd7, 1'd1} : pll_fbdiv_ring_fbck_expected = 10'b0000100000;
default: pll_fbdiv_ring_fbck_expected = 10'bzzzzzzzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel} )
  {PCIE, 4'd0, 5'd0, 1'd0} : icp_ring_expected = 4'b1111;
  {PCIE, 4'd0, 5'd1, 1'd0} : icp_ring_expected = 4'b1101;
  {PCIE, 4'd0, 5'd2, 1'd0} : icp_ring_expected = 4'b1101;
  {PCIE, 4'd0, 5'd3, 1'd0} : icp_ring_expected = 4'b1100;
  {PCIE, 4'd0, 5'd4, 1'd0} : icp_ring_expected = 4'b1100;
  {PCIE, 4'd0, 5'd5, 1'd0} : icp_ring_expected = 4'b1111;
  {PCIE, 4'd0, 5'd6, 1'd0} : icp_ring_expected = 4'b1101;
  {PCIE, 4'd0, 5'd7, 1'd0} : icp_ring_expected = 4'b1101;
  {PCIE, 4'd1, 5'd0, 1'd0} : icp_ring_expected = 4'b1111;
  {PCIE, 4'd1, 5'd1, 1'd0} : icp_ring_expected = 4'b1101;
  {PCIE, 4'd1, 5'd2, 1'd0} : icp_ring_expected = 4'b1101;
  {PCIE, 4'd1, 5'd3, 1'd0} : icp_ring_expected = 4'b1100;
  {PCIE, 4'd1, 5'd4, 1'd0} : icp_ring_expected = 4'b1100;
  {PCIE, 4'd1, 5'd5, 1'd0} : icp_ring_expected = 4'b1111;
  {PCIE, 4'd1, 5'd6, 1'd0} : icp_ring_expected = 4'b1101;
  {PCIE, 4'd1, 5'd7, 1'd0} : icp_ring_expected = 4'b1101;
  {PCIE, 4'd0, 5'd0, 1'd1} : icp_ring_expected = 4'b1111;
  {PCIE, 4'd0, 5'd1, 1'd1} : icp_ring_expected = 4'b1110;
  {PCIE, 4'd0, 5'd2, 1'd1} : icp_ring_expected = 4'b1100;
  {PCIE, 4'd0, 5'd3, 1'd1} : icp_ring_expected = 4'b1101;
  {PCIE, 4'd0, 5'd4, 1'd1} : icp_ring_expected = 4'b1100;
  {PCIE, 4'd0, 5'd5, 1'd1} : icp_ring_expected = 4'b1111;
  {PCIE, 4'd0, 5'd6, 1'd1} : icp_ring_expected = 4'b1101;
  {PCIE, 4'd0, 5'd7, 1'd1} : icp_ring_expected = 4'b1111;
  {PCIE, 4'd1, 5'd0, 1'd1} : icp_ring_expected = 4'b1111;
  {PCIE, 4'd1, 5'd1, 1'd1} : icp_ring_expected = 4'b1110;
  {PCIE, 4'd1, 5'd2, 1'd1} : icp_ring_expected = 4'b1100;
  {PCIE, 4'd1, 5'd3, 1'd1} : icp_ring_expected = 4'b1101;
  {PCIE, 4'd1, 5'd4, 1'd1} : icp_ring_expected = 4'b1100;
  {PCIE, 4'd1, 5'd5, 1'd1} : icp_ring_expected = 4'b1111;
  {PCIE, 4'd1, 5'd6, 1'd1} : icp_ring_expected = 4'b1101;
  {PCIE, 4'd1, 5'd7, 1'd1} : icp_ring_expected = 4'b1111;
default: icp_ring_expected = 4'bzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel} )
  {PCIE, 4'd0, 5'd0, 1'd0} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd0, 5'd1, 1'd0} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd0, 5'd2, 1'd0} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd0, 5'd3, 1'd0} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd0, 5'd4, 1'd0} : pll_speed_thresh_ring_expected = 9'b011111100;
  {PCIE, 4'd0, 5'd5, 1'd0} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd0, 5'd6, 1'd0} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd0, 5'd7, 1'd0} : pll_speed_thresh_ring_expected = 9'b011111011;
  {PCIE, 4'd1, 5'd0, 1'd0} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd1, 5'd1, 1'd0} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd1, 5'd2, 1'd0} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd1, 5'd3, 1'd0} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd1, 5'd4, 1'd0} : pll_speed_thresh_ring_expected = 9'b011111100;
  {PCIE, 4'd1, 5'd5, 1'd0} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd1, 5'd6, 1'd0} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd1, 5'd7, 1'd0} : pll_speed_thresh_ring_expected = 9'b011111011;
  {PCIE, 4'd0, 5'd0, 1'd1} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd0, 5'd1, 1'd1} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd0, 5'd2, 1'd1} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd0, 5'd3, 1'd1} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd0, 5'd4, 1'd1} : pll_speed_thresh_ring_expected = 9'b011111100;
  {PCIE, 4'd0, 5'd5, 1'd1} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd0, 5'd6, 1'd1} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd0, 5'd7, 1'd1} : pll_speed_thresh_ring_expected = 9'b011111011;
  {PCIE, 4'd1, 5'd0, 1'd1} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd1, 5'd1, 1'd1} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd1, 5'd2, 1'd1} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd1, 5'd3, 1'd1} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd1, 5'd4, 1'd1} : pll_speed_thresh_ring_expected = 9'b011111100;
  {PCIE, 4'd1, 5'd5, 1'd1} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd1, 5'd6, 1'd1} : pll_speed_thresh_ring_expected = 9'b011111010;
  {PCIE, 4'd1, 5'd7, 1'd1} : pll_speed_thresh_ring_expected = 9'b011111011;
default: pll_speed_thresh_ring_expected = 9'bzzzzzzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel} )
  {PCIE, 4'd0, 5'd0, 1'd0} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd0, 5'd1, 1'd0} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd0, 5'd2, 1'd0} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd0, 5'd3, 1'd0} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd0, 5'd4, 1'd0} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd0, 5'd5, 1'd0} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd0, 5'd6, 1'd0} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd0, 5'd7, 1'd0} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd1, 5'd0, 1'd0} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd1, 5'd1, 1'd0} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd1, 5'd2, 1'd0} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd1, 5'd3, 1'd0} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd1, 5'd4, 1'd0} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd1, 5'd5, 1'd0} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd1, 5'd6, 1'd0} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd1, 5'd7, 1'd0} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd0, 5'd0, 1'd1} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd0, 5'd1, 1'd1} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd0, 5'd2, 1'd1} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd0, 5'd3, 1'd1} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd0, 5'd4, 1'd1} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd0, 5'd5, 1'd1} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd0, 5'd6, 1'd1} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd0, 5'd7, 1'd1} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd1, 5'd0, 1'd1} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd1, 5'd1, 1'd1} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd1, 5'd2, 1'd1} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd1, 5'd3, 1'd1} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd1, 5'd4, 1'd1} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd1, 5'd5, 1'd1} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd1, 5'd6, 1'd1} : fbdiv_cal_ring_expected = 10'b0000101000;
  {PCIE, 4'd1, 5'd7, 1'd1} : fbdiv_cal_ring_expected = 10'b0000101000;
default: fbdiv_cal_ring_expected = 10'bzzzzzzzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel} )
  {PCIE, 4'd0, 5'd0, 1'd0} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd0, 5'd1, 1'd0} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd0, 5'd2, 1'd0} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd0, 5'd3, 1'd0} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd0, 5'd4, 1'd0} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd0, 5'd5, 1'd0} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd0, 5'd6, 1'd0} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd0, 5'd7, 1'd0} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd1, 5'd0, 1'd0} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd1, 5'd1, 1'd0} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd1, 5'd2, 1'd0} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd1, 5'd3, 1'd0} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd1, 5'd4, 1'd0} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd1, 5'd5, 1'd0} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd1, 5'd6, 1'd0} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd1, 5'd7, 1'd0} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd0, 5'd0, 1'd1} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd0, 5'd1, 1'd1} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd0, 5'd2, 1'd1} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd0, 5'd3, 1'd1} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd0, 5'd4, 1'd1} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd0, 5'd5, 1'd1} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd0, 5'd6, 1'd1} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd0, 5'd7, 1'd1} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd1, 5'd0, 1'd1} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd1, 5'd1, 1'd1} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd1, 5'd2, 1'd1} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd1, 5'd3, 1'd1} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd1, 5'd4, 1'd1} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd1, 5'd5, 1'd1} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd1, 5'd6, 1'd1} : intpi_ring_expected = 4'b0101;
  {PCIE, 4'd1, 5'd7, 1'd1} : intpi_ring_expected = 4'b0101;
default: intpi_ring_expected = 4'bzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel} )
  {PCIE, 4'd0, 5'd0, 1'd0} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd0, 5'd1, 1'd0} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd0, 5'd2, 1'd0} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd0, 5'd3, 1'd0} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd0, 5'd4, 1'd0} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd0, 5'd5, 1'd0} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd0, 5'd6, 1'd0} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd0, 5'd7, 1'd0} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd1, 5'd0, 1'd0} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd1, 5'd1, 1'd0} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd1, 5'd2, 1'd0} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd1, 5'd3, 1'd0} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd1, 5'd4, 1'd0} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd1, 5'd5, 1'd0} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd1, 5'd6, 1'd0} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd1, 5'd7, 1'd0} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd0, 5'd0, 1'd1} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd0, 5'd1, 1'd1} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd0, 5'd2, 1'd1} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd0, 5'd3, 1'd1} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd0, 5'd4, 1'd1} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd0, 5'd5, 1'd1} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd0, 5'd6, 1'd1} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd0, 5'd7, 1'd1} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd1, 5'd0, 1'd1} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd1, 5'd1, 1'd1} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd1, 5'd2, 1'd1} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd1, 5'd3, 1'd1} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd1, 5'd4, 1'd1} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd1, 5'd5, 1'd1} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd1, 5'd6, 1'd1} : tx_intpr_ring_expected = 2'b10;
  {PCIE, 4'd1, 5'd7, 1'd1} : tx_intpr_ring_expected = 2'b10;
default: tx_intpr_ring_expected = 2'bzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel} )
  {PCIE, 4'd0, 5'd0, 1'd0} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd1, 1'd0} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd2, 1'd0} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd3, 1'd0} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd4, 1'd0} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd5, 1'd0} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd6, 1'd0} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd7, 1'd0} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd0, 1'd0} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd1, 1'd0} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd2, 1'd0} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd3, 1'd0} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd4, 1'd0} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd5, 1'd0} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd6, 1'd0} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd7, 1'd0} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd0, 1'd1} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd1, 1'd1} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd2, 1'd1} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd3, 1'd1} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd4, 1'd1} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd5, 1'd1} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd6, 1'd1} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd7, 1'd1} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd0, 1'd1} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd1, 1'd1} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd2, 1'd1} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd3, 1'd1} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd4, 1'd1} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd5, 1'd1} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd6, 1'd1} : pll_band_sel_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd7, 1'd1} : pll_band_sel_ring_expected = 1'b0;
default: pll_band_sel_ring_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel} )
  {PCIE, 4'd0, 5'd0, 1'd0} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd0, 5'd1, 1'd0} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd0, 5'd2, 1'd0} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd0, 5'd3, 1'd0} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd0, 5'd4, 1'd0} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd0, 5'd5, 1'd0} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd0, 5'd6, 1'd0} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd0, 5'd7, 1'd0} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd1, 5'd0, 1'd0} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd1, 5'd1, 1'd0} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd1, 5'd2, 1'd0} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd1, 5'd3, 1'd0} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd1, 5'd4, 1'd0} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd1, 5'd5, 1'd0} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd1, 5'd6, 1'd0} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd1, 5'd7, 1'd0} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd0, 5'd0, 1'd1} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd0, 5'd1, 1'd1} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd0, 5'd2, 1'd1} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd0, 5'd3, 1'd1} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd0, 5'd4, 1'd1} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd0, 5'd5, 1'd1} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd0, 5'd6, 1'd1} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd0, 5'd7, 1'd1} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd1, 5'd0, 1'd1} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd1, 5'd1, 1'd1} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd1, 5'd2, 1'd1} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd1, 5'd3, 1'd1} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd1, 5'd4, 1'd1} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd1, 5'd5, 1'd1} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd1, 5'd6, 1'd1} : pll_lpf_c1_sel_ring_expected = 2'b11;
  {PCIE, 4'd1, 5'd7, 1'd1} : pll_lpf_c1_sel_ring_expected = 2'b11;
default: pll_lpf_c1_sel_ring_expected = 2'bzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel} )
  {PCIE, 4'd0, 5'd0, 1'd0} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd0, 5'd1, 1'd0} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd0, 5'd2, 1'd0} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd0, 5'd3, 1'd0} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd0, 5'd4, 1'd0} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd0, 5'd5, 1'd0} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd0, 5'd6, 1'd0} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd0, 5'd7, 1'd0} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd1, 5'd0, 1'd0} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd1, 5'd1, 1'd0} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd1, 5'd2, 1'd0} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd1, 5'd3, 1'd0} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd1, 5'd4, 1'd0} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd1, 5'd5, 1'd0} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd1, 5'd6, 1'd0} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd1, 5'd7, 1'd0} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd0, 5'd0, 1'd1} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd0, 5'd1, 1'd1} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd0, 5'd2, 1'd1} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd0, 5'd3, 1'd1} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd0, 5'd4, 1'd1} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd0, 5'd5, 1'd1} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd0, 5'd6, 1'd1} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd0, 5'd7, 1'd1} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd1, 5'd0, 1'd1} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd1, 5'd1, 1'd1} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd1, 5'd2, 1'd1} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd1, 5'd3, 1'd1} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd1, 5'd4, 1'd1} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd1, 5'd5, 1'd1} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd1, 5'd6, 1'd1} : pll_lpf_c2_sel_ring_expected = 2'b00;
  {PCIE, 4'd1, 5'd7, 1'd1} : pll_lpf_c2_sel_ring_expected = 2'b00;
default: pll_lpf_c2_sel_ring_expected = 2'bzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel} )
  {PCIE, 4'd0, 5'd0, 1'd0} : pll_lpf_r1_sel_ring_expected = 3'b001;
  {PCIE, 4'd0, 5'd1, 1'd0} : pll_lpf_r1_sel_ring_expected = 3'b001;
  {PCIE, 4'd0, 5'd2, 1'd0} : pll_lpf_r1_sel_ring_expected = 3'b001;
  {PCIE, 4'd0, 5'd3, 1'd0} : pll_lpf_r1_sel_ring_expected = 3'b010;
  {PCIE, 4'd0, 5'd4, 1'd0} : pll_lpf_r1_sel_ring_expected = 3'b010;
  {PCIE, 4'd0, 5'd5, 1'd0} : pll_lpf_r1_sel_ring_expected = 3'b001;
  {PCIE, 4'd0, 5'd6, 1'd0} : pll_lpf_r1_sel_ring_expected = 3'b100;
  {PCIE, 4'd0, 5'd7, 1'd0} : pll_lpf_r1_sel_ring_expected = 3'b101;
  {PCIE, 4'd1, 5'd0, 1'd0} : pll_lpf_r1_sel_ring_expected = 3'b001;
  {PCIE, 4'd1, 5'd1, 1'd0} : pll_lpf_r1_sel_ring_expected = 3'b001;
  {PCIE, 4'd1, 5'd2, 1'd0} : pll_lpf_r1_sel_ring_expected = 3'b001;
  {PCIE, 4'd1, 5'd3, 1'd0} : pll_lpf_r1_sel_ring_expected = 3'b010;
  {PCIE, 4'd1, 5'd4, 1'd0} : pll_lpf_r1_sel_ring_expected = 3'b010;
  {PCIE, 4'd1, 5'd5, 1'd0} : pll_lpf_r1_sel_ring_expected = 3'b001;
  {PCIE, 4'd1, 5'd6, 1'd0} : pll_lpf_r1_sel_ring_expected = 3'b100;
  {PCIE, 4'd1, 5'd7, 1'd0} : pll_lpf_r1_sel_ring_expected = 3'b101;
  {PCIE, 4'd0, 5'd0, 1'd1} : pll_lpf_r1_sel_ring_expected = 3'b001;
  {PCIE, 4'd0, 5'd1, 1'd1} : pll_lpf_r1_sel_ring_expected = 3'b001;
  {PCIE, 4'd0, 5'd2, 1'd1} : pll_lpf_r1_sel_ring_expected = 3'b001;
  {PCIE, 4'd0, 5'd3, 1'd1} : pll_lpf_r1_sel_ring_expected = 3'b010;
  {PCIE, 4'd0, 5'd4, 1'd1} : pll_lpf_r1_sel_ring_expected = 3'b010;
  {PCIE, 4'd0, 5'd5, 1'd1} : pll_lpf_r1_sel_ring_expected = 3'b001;
  {PCIE, 4'd0, 5'd6, 1'd1} : pll_lpf_r1_sel_ring_expected = 3'b100;
  {PCIE, 4'd0, 5'd7, 1'd1} : pll_lpf_r1_sel_ring_expected = 3'b100;
  {PCIE, 4'd1, 5'd0, 1'd1} : pll_lpf_r1_sel_ring_expected = 3'b001;
  {PCIE, 4'd1, 5'd1, 1'd1} : pll_lpf_r1_sel_ring_expected = 3'b001;
  {PCIE, 4'd1, 5'd2, 1'd1} : pll_lpf_r1_sel_ring_expected = 3'b001;
  {PCIE, 4'd1, 5'd3, 1'd1} : pll_lpf_r1_sel_ring_expected = 3'b010;
  {PCIE, 4'd1, 5'd4, 1'd1} : pll_lpf_r1_sel_ring_expected = 3'b010;
  {PCIE, 4'd1, 5'd5, 1'd1} : pll_lpf_r1_sel_ring_expected = 3'b001;
  {PCIE, 4'd1, 5'd6, 1'd1} : pll_lpf_r1_sel_ring_expected = 3'b100;
  {PCIE, 4'd1, 5'd7, 1'd1} : pll_lpf_r1_sel_ring_expected = 3'b100;
default: pll_lpf_r1_sel_ring_expected = 3'bzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel} )
  {PCIE, 4'd0, 5'd0, 1'd0} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd1, 1'd0} : init_txfoffs_ring_expected = 10'b1111011111;
  {PCIE, 4'd0, 5'd2, 1'd0} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd3, 1'd0} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd4, 1'd0} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd5, 1'd0} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd6, 1'd0} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd7, 1'd0} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd0, 1'd0} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd1, 1'd0} : init_txfoffs_ring_expected = 10'b1111011111;
  {PCIE, 4'd1, 5'd2, 1'd0} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd3, 1'd0} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd4, 1'd0} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd5, 1'd0} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd6, 1'd0} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd7, 1'd0} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd0, 1'd1} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd1, 1'd1} : init_txfoffs_ring_expected = 10'b1101111101;
  {PCIE, 4'd0, 5'd2, 1'd1} : init_txfoffs_ring_expected = 10'b1011111010;
  {PCIE, 4'd0, 5'd3, 1'd1} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd4, 1'd1} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd5, 1'd1} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd6, 1'd1} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd7, 1'd1} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd0, 1'd1} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd1, 1'd1} : init_txfoffs_ring_expected = 10'b1101111101;
  {PCIE, 4'd1, 5'd2, 1'd1} : init_txfoffs_ring_expected = 10'b1011111010;
  {PCIE, 4'd1, 5'd3, 1'd1} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd4, 1'd1} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd5, 1'd1} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd6, 1'd1} : init_txfoffs_ring_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd7, 1'd1} : init_txfoffs_ring_expected = 10'b0000000000;
default: init_txfoffs_ring_expected = 10'bzzzzzzzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel} )
  {PCIE, 4'd0, 5'd0, 1'd0} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd1, 1'd0} : init_txfoffs_ring_fbck_expected = 10'b1111011111;
  {PCIE, 4'd0, 5'd2, 1'd0} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd3, 1'd0} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd4, 1'd0} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd5, 1'd0} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd6, 1'd0} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd7, 1'd0} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd0, 1'd0} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd1, 1'd0} : init_txfoffs_ring_fbck_expected = 10'b1111011111;
  {PCIE, 4'd1, 5'd2, 1'd0} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd3, 1'd0} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd4, 1'd0} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd5, 1'd0} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd6, 1'd0} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd7, 1'd0} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd0, 1'd1} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd1, 1'd1} : init_txfoffs_ring_fbck_expected = 10'b1101111101;
  {PCIE, 4'd0, 5'd2, 1'd1} : init_txfoffs_ring_fbck_expected = 10'b1011111010;
  {PCIE, 4'd0, 5'd3, 1'd1} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd4, 1'd1} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd5, 1'd1} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd6, 1'd1} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd0, 5'd7, 1'd1} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd0, 1'd1} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd1, 1'd1} : init_txfoffs_ring_fbck_expected = 10'b1101111101;
  {PCIE, 4'd1, 5'd2, 1'd1} : init_txfoffs_ring_fbck_expected = 10'b1011111010;
  {PCIE, 4'd1, 5'd3, 1'd1} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd4, 1'd1} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd5, 1'd1} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd6, 1'd1} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
  {PCIE, 4'd1, 5'd7, 1'd1} : init_txfoffs_ring_fbck_expected = 10'b0000000000;
default: init_txfoffs_ring_fbck_expected = 10'bzzzzzzzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel} )
  {PCIE, 4'd0, 5'd0, 1'd0} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd1, 1'd0} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd2, 1'd0} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd3, 1'd0} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd4, 1'd0} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd5, 1'd0} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd6, 1'd0} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd7, 1'd0} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd0, 1'd0} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd1, 1'd0} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd2, 1'd0} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd3, 1'd0} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd4, 1'd0} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd5, 1'd0} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd6, 1'd0} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd7, 1'd0} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd0, 1'd1} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd1, 1'd1} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd2, 1'd1} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd3, 1'd1} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd4, 1'd1} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd5, 1'd1} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd6, 1'd1} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd0, 5'd7, 1'd1} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd0, 1'd1} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd1, 1'd1} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd2, 1'd1} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd3, 1'd1} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd4, 1'd1} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd5, 1'd1} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd6, 1'd1} : ssc_acc_factor_ring_expected = 1'b0;
  {PCIE, 4'd1, 5'd7, 1'd1} : ssc_acc_factor_ring_expected = 1'b0;
default: ssc_acc_factor_ring_expected = 1'bz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel} )
  {PCIE, 4'd0, 5'd0, 1'd0} : ssc_step_125ppm_ring_expected = 4'b0000;
  {PCIE, 4'd0, 5'd1, 1'd0} : ssc_step_125ppm_ring_expected = 4'b0000;
  {PCIE, 4'd0, 5'd2, 1'd0} : ssc_step_125ppm_ring_expected = 4'b0000;
  {PCIE, 4'd0, 5'd3, 1'd0} : ssc_step_125ppm_ring_expected = 4'b0000;
  {PCIE, 4'd0, 5'd4, 1'd0} : ssc_step_125ppm_ring_expected = 4'b0000;
  {PCIE, 4'd0, 5'd5, 1'd0} : ssc_step_125ppm_ring_expected = 4'b0000;
  {PCIE, 4'd0, 5'd6, 1'd0} : ssc_step_125ppm_ring_expected = 4'b0000;
  {PCIE, 4'd0, 5'd7, 1'd0} : ssc_step_125ppm_ring_expected = 4'b0000;
  {PCIE, 4'd1, 5'd0, 1'd0} : ssc_step_125ppm_ring_expected = 4'b0000;
  {PCIE, 4'd1, 5'd1, 1'd0} : ssc_step_125ppm_ring_expected = 4'b0000;
  {PCIE, 4'd1, 5'd2, 1'd0} : ssc_step_125ppm_ring_expected = 4'b0000;
  {PCIE, 4'd1, 5'd3, 1'd0} : ssc_step_125ppm_ring_expected = 4'b0000;
  {PCIE, 4'd1, 5'd4, 1'd0} : ssc_step_125ppm_ring_expected = 4'b0000;
  {PCIE, 4'd1, 5'd5, 1'd0} : ssc_step_125ppm_ring_expected = 4'b0000;
  {PCIE, 4'd1, 5'd6, 1'd0} : ssc_step_125ppm_ring_expected = 4'b0000;
  {PCIE, 4'd1, 5'd7, 1'd0} : ssc_step_125ppm_ring_expected = 4'b0000;
  {PCIE, 4'd0, 5'd0, 1'd1} : ssc_step_125ppm_ring_expected = 4'b0011;
  {PCIE, 4'd0, 5'd1, 1'd1} : ssc_step_125ppm_ring_expected = 4'b0011;
  {PCIE, 4'd0, 5'd2, 1'd1} : ssc_step_125ppm_ring_expected = 4'b0011;
  {PCIE, 4'd0, 5'd3, 1'd1} : ssc_step_125ppm_ring_expected = 4'b0011;
  {PCIE, 4'd0, 5'd4, 1'd1} : ssc_step_125ppm_ring_expected = 4'b0011;
  {PCIE, 4'd0, 5'd5, 1'd1} : ssc_step_125ppm_ring_expected = 4'b0011;
  {PCIE, 4'd0, 5'd6, 1'd1} : ssc_step_125ppm_ring_expected = 4'b0011;
  {PCIE, 4'd0, 5'd7, 1'd1} : ssc_step_125ppm_ring_expected = 4'b0011;
  {PCIE, 4'd1, 5'd0, 1'd1} : ssc_step_125ppm_ring_expected = 4'b0011;
  {PCIE, 4'd1, 5'd1, 1'd1} : ssc_step_125ppm_ring_expected = 4'b0011;
  {PCIE, 4'd1, 5'd2, 1'd1} : ssc_step_125ppm_ring_expected = 4'b0011;
  {PCIE, 4'd1, 5'd3, 1'd1} : ssc_step_125ppm_ring_expected = 4'b0011;
  {PCIE, 4'd1, 5'd4, 1'd1} : ssc_step_125ppm_ring_expected = 4'b0011;
  {PCIE, 4'd1, 5'd5, 1'd1} : ssc_step_125ppm_ring_expected = 4'b0011;
  {PCIE, 4'd1, 5'd6, 1'd1} : ssc_step_125ppm_ring_expected = 4'b0011;
  {PCIE, 4'd1, 5'd7, 1'd1} : ssc_step_125ppm_ring_expected = 4'b0011;
default: ssc_step_125ppm_ring_expected = 4'bzzzz;

endcase

always @(phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel)
case ( {phy_mode_bit[2:0], gen[3:0], refclk_fsel_ring[4:0], reg_fbck_sel} )
  {PCIE, 4'd0, 5'd0, 1'd0} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd0, 5'd1, 1'd0} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd0, 5'd2, 1'd0} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd0, 5'd3, 1'd0} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd0, 5'd4, 1'd0} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd0, 5'd5, 1'd0} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd0, 5'd6, 1'd0} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd0, 5'd7, 1'd0} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd1, 5'd0, 1'd0} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd1, 5'd1, 1'd0} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd1, 5'd2, 1'd0} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd1, 5'd3, 1'd0} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd1, 5'd4, 1'd0} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd1, 5'd5, 1'd0} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd1, 5'd6, 1'd0} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd1, 5'd7, 1'd0} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd0, 5'd0, 1'd1} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd0, 5'd1, 1'd1} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd0, 5'd2, 1'd1} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd0, 5'd3, 1'd1} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd0, 5'd4, 1'd1} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd0, 5'd5, 1'd1} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd0, 5'd6, 1'd1} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd0, 5'd7, 1'd1} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd1, 5'd0, 1'd1} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd1, 5'd1, 1'd1} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd1, 5'd2, 1'd1} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd1, 5'd3, 1'd1} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd1, 5'd4, 1'd1} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd1, 5'd5, 1'd1} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd1, 5'd6, 1'd1} : ssc_m_ring_expected = 13'b0100110101111;
  {PCIE, 4'd1, 5'd7, 1'd1} : ssc_m_ring_expected = 13'b0100110101111;
default: ssc_m_ring_expected = 13'bzzzzzzzzzzzzz;

endcase


endmodule
`endif